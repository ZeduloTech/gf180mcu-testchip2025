VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_wb_mem_64x32
  CLASS BLOCK ;
  FOREIGN efuse_wb_mem_64x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 204.530 BY 1311.065 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.080 2.760 6.080 1306.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 2.760 200.320 4.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 1304.520 200.320 1306.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.320 2.760 200.320 1306.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 0.260 15.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 1286.625 15.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.280 0.260 65.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 0.260 115.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 1285.580 115.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 0.260 165.880 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 15.960 202.820 17.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 65.960 202.820 67.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 115.960 202.820 117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 165.960 202.820 167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 215.960 202.820 217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 265.960 202.820 267.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 315.960 202.820 317.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 365.960 202.820 367.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 415.960 202.820 417.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 465.960 202.820 467.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 515.960 202.820 517.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 565.960 202.820 567.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 615.960 202.820 617.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 665.960 202.820 667.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 715.960 202.820 717.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 765.960 202.820 767.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 815.960 202.820 817.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 865.960 202.820 867.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 915.960 202.820 917.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 965.960 202.820 967.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1015.960 202.820 1017.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1065.960 202.820 1067.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1115.960 202.820 1117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1165.960 202.820 1167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1215.960 202.820 1217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1265.960 202.820 1267.560 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 1.580 0.260 3.580 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 0.260 202.820 2.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1307.020 202.820 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.820 0.260 202.820 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 0.260 19.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 1286.000 19.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.580 0.260 69.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 0.260 119.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 1286.000 119.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 0.260 169.180 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 19.260 202.820 20.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 69.260 202.820 70.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 119.260 202.820 120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 169.260 202.820 170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 219.260 202.820 220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 269.260 202.820 270.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 319.260 202.820 320.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 369.260 202.820 370.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 419.260 202.820 420.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 469.260 202.820 470.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 519.260 202.820 520.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 569.260 202.820 570.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 619.260 202.820 620.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 669.260 202.820 670.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 719.260 202.820 720.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 769.260 202.820 770.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 819.260 202.820 820.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 869.260 202.820 870.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 919.260 202.820 920.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 969.260 202.820 970.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1019.260 202.820 1020.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1069.260 202.820 1070.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1119.260 202.820 1120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1169.260 202.820 1170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1219.260 202.820 1220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1269.260 202.820 1270.860 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1310.505 17.360 1311.065 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 1310.505 26.320 1311.065 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 1310.505 28.560 1311.065 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 1310.505 30.800 1311.065 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 1310.505 33.040 1311.065 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 1310.505 35.280 1311.065 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 1310.505 37.520 1311.065 ;
    END
  END wb_adr_i[5]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 1310.505 21.840 1311.065 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 1310.505 15.120 1311.065 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 1310.505 39.760 1311.065 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 1310.505 62.160 1311.065 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 1310.505 64.400 1311.065 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 1310.505 66.640 1311.065 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 1310.505 68.880 1311.065 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1310.505 71.120 1311.065 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 1310.505 73.360 1311.065 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 1310.505 75.600 1311.065 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1310.505 77.840 1311.065 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 1310.505 80.080 1311.065 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 1310.505 82.320 1311.065 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 1310.505 42.000 1311.065 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1310.505 84.560 1311.065 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 1310.505 86.800 1311.065 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 1310.505 89.040 1311.065 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1310.505 91.280 1311.065 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 1310.505 93.520 1311.065 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 1310.505 95.760 1311.065 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1310.505 98.000 1311.065 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 1310.505 100.240 1311.065 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 1310.505 102.480 1311.065 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1310.505 104.720 1311.065 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1310.505 44.240 1311.065 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 1310.505 106.960 1311.065 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 1310.505 109.200 1311.065 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 1310.505 46.480 1311.065 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 1310.505 48.720 1311.065 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1310.505 50.960 1311.065 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 1310.505 53.200 1311.065 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 1310.505 55.440 1311.065 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1310.505 57.680 1311.065 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 1310.505 59.920 1311.065 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 1310.505 120.400 1311.065 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 1310.505 142.800 1311.065 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1310.505 145.040 1311.065 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 1310.505 147.280 1311.065 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 1310.505 149.520 1311.065 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1310.505 151.760 1311.065 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 1310.505 154.000 1311.065 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 1310.505 156.240 1311.065 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1310.505 158.480 1311.065 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 1310.505 160.720 1311.065 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 1310.505 162.960 1311.065 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 1310.505 122.640 1311.065 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 1310.505 165.200 1311.065 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 1310.505 167.440 1311.065 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 1310.505 169.680 1311.065 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1310.505 171.920 1311.065 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 1310.505 174.160 1311.065 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 1310.505 176.400 1311.065 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1310.505 178.640 1311.065 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 1310.505 180.880 1311.065 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 1310.505 183.120 1311.065 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1310.505 185.360 1311.065 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1310.505 124.880 1311.065 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 1310.505 187.600 1311.065 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 1310.505 189.840 1311.065 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 1310.505 127.120 1311.065 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 1310.505 129.360 1311.065 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 1310.505 131.600 1311.065 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 1310.505 133.840 1311.065 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 1310.505 136.080 1311.065 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 1310.505 138.320 1311.065 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 1310.505 140.560 1311.065 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 1310.505 19.600 1311.065 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1310.505 111.440 1311.065 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 1310.505 113.680 1311.065 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 1310.505 115.920 1311.065 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 1310.505 118.160 1311.065 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 1310.505 12.880 1311.065 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1310.505 24.080 1311.065 ;
    END
  END wb_we_i
  PIN write_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.528000 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1310.505 192.080 1311.065 ;
    END
  END write_enable_i
  OBS
      LAYER Nwell ;
        RECT 9.650 11.330 194.750 1297.950 ;
      LAYER Metal1 ;
        RECT 10.080 11.460 194.320 1297.820 ;
      LAYER Metal2 ;
        RECT 0.140 1310.205 12.020 1310.505 ;
        RECT 13.180 1310.205 14.260 1310.505 ;
        RECT 15.420 1310.205 16.500 1310.505 ;
        RECT 17.660 1310.205 18.740 1310.505 ;
        RECT 19.900 1310.205 20.980 1310.505 ;
        RECT 22.140 1310.205 23.220 1310.505 ;
        RECT 24.380 1310.205 25.460 1310.505 ;
        RECT 26.620 1310.205 27.700 1310.505 ;
        RECT 28.860 1310.205 29.940 1310.505 ;
        RECT 31.100 1310.205 32.180 1310.505 ;
        RECT 33.340 1310.205 34.420 1310.505 ;
        RECT 35.580 1310.205 36.660 1310.505 ;
        RECT 37.820 1310.205 38.900 1310.505 ;
        RECT 40.060 1310.205 41.140 1310.505 ;
        RECT 42.300 1310.205 43.380 1310.505 ;
        RECT 44.540 1310.205 45.620 1310.505 ;
        RECT 46.780 1310.205 47.860 1310.505 ;
        RECT 49.020 1310.205 50.100 1310.505 ;
        RECT 51.260 1310.205 52.340 1310.505 ;
        RECT 53.500 1310.205 54.580 1310.505 ;
        RECT 55.740 1310.205 56.820 1310.505 ;
        RECT 57.980 1310.205 59.060 1310.505 ;
        RECT 60.220 1310.205 61.300 1310.505 ;
        RECT 62.460 1310.205 63.540 1310.505 ;
        RECT 64.700 1310.205 65.780 1310.505 ;
        RECT 66.940 1310.205 68.020 1310.505 ;
        RECT 69.180 1310.205 70.260 1310.505 ;
        RECT 71.420 1310.205 72.500 1310.505 ;
        RECT 73.660 1310.205 74.740 1310.505 ;
        RECT 75.900 1310.205 76.980 1310.505 ;
        RECT 78.140 1310.205 79.220 1310.505 ;
        RECT 80.380 1310.205 81.460 1310.505 ;
        RECT 82.620 1310.205 83.700 1310.505 ;
        RECT 84.860 1310.205 85.940 1310.505 ;
        RECT 87.100 1310.205 88.180 1310.505 ;
        RECT 89.340 1310.205 90.420 1310.505 ;
        RECT 91.580 1310.205 92.660 1310.505 ;
        RECT 93.820 1310.205 94.900 1310.505 ;
        RECT 96.060 1310.205 97.140 1310.505 ;
        RECT 98.300 1310.205 99.380 1310.505 ;
        RECT 100.540 1310.205 101.620 1310.505 ;
        RECT 102.780 1310.205 103.860 1310.505 ;
        RECT 105.020 1310.205 106.100 1310.505 ;
        RECT 107.260 1310.205 108.340 1310.505 ;
        RECT 109.500 1310.205 110.580 1310.505 ;
        RECT 111.740 1310.205 112.820 1310.505 ;
        RECT 113.980 1310.205 115.060 1310.505 ;
        RECT 116.220 1310.205 117.300 1310.505 ;
        RECT 118.460 1310.205 119.540 1310.505 ;
        RECT 120.700 1310.205 121.780 1310.505 ;
        RECT 122.940 1310.205 124.020 1310.505 ;
        RECT 125.180 1310.205 126.260 1310.505 ;
        RECT 127.420 1310.205 128.500 1310.505 ;
        RECT 129.660 1310.205 130.740 1310.505 ;
        RECT 131.900 1310.205 132.980 1310.505 ;
        RECT 134.140 1310.205 135.220 1310.505 ;
        RECT 136.380 1310.205 137.460 1310.505 ;
        RECT 138.620 1310.205 139.700 1310.505 ;
        RECT 140.860 1310.205 141.940 1310.505 ;
        RECT 143.100 1310.205 144.180 1310.505 ;
        RECT 145.340 1310.205 146.420 1310.505 ;
        RECT 147.580 1310.205 148.660 1310.505 ;
        RECT 149.820 1310.205 150.900 1310.505 ;
        RECT 152.060 1310.205 153.140 1310.505 ;
        RECT 154.300 1310.205 155.380 1310.505 ;
        RECT 156.540 1310.205 157.620 1310.505 ;
        RECT 158.780 1310.205 159.860 1310.505 ;
        RECT 161.020 1310.205 162.100 1310.505 ;
        RECT 163.260 1310.205 164.340 1310.505 ;
        RECT 165.500 1310.205 166.580 1310.505 ;
        RECT 167.740 1310.205 168.820 1310.505 ;
        RECT 169.980 1310.205 171.060 1310.505 ;
        RECT 172.220 1310.205 173.300 1310.505 ;
        RECT 174.460 1310.205 175.540 1310.505 ;
        RECT 176.700 1310.205 177.780 1310.505 ;
        RECT 178.940 1310.205 180.020 1310.505 ;
        RECT 181.180 1310.205 182.260 1310.505 ;
        RECT 183.420 1310.205 184.500 1310.505 ;
        RECT 185.660 1310.205 186.740 1310.505 ;
        RECT 187.900 1310.205 188.980 1310.505 ;
        RECT 190.140 1310.205 191.220 1310.505 ;
        RECT 192.380 1310.205 204.260 1310.505 ;
        RECT 0.140 11.570 204.260 1310.205 ;
      LAYER Metal3 ;
        RECT 0.090 7.420 204.310 1310.260 ;
      LAYER Metal4 ;
        RECT 0.140 1309.320 204.260 1310.310 ;
        RECT 0.140 7.370 1.280 1309.320 ;
        RECT 3.880 1306.820 13.980 1309.320 ;
        RECT 6.380 1286.325 13.980 1306.820 ;
        RECT 16.180 1286.325 17.280 1309.320 ;
        RECT 6.380 1285.700 17.280 1286.325 ;
        RECT 19.480 1285.700 63.980 1309.320 ;
        RECT 6.380 7.370 63.980 1285.700 ;
        RECT 66.180 7.370 67.280 1309.320 ;
        RECT 69.480 1285.280 113.980 1309.320 ;
        RECT 116.180 1285.700 117.280 1309.320 ;
        RECT 119.480 1285.700 163.980 1309.320 ;
        RECT 116.180 1285.280 163.980 1285.700 ;
        RECT 69.480 7.370 163.980 1285.280 ;
        RECT 166.180 7.370 167.280 1309.320 ;
        RECT 169.480 1306.820 200.520 1309.320 ;
        RECT 169.480 7.370 198.020 1306.820 ;
        RECT 203.120 7.370 204.260 1309.320 ;
  END
END efuse_wb_mem_64x32
END LIBRARY

