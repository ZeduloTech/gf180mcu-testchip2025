module efuse_wb_mem_64x32 (wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rst_i,
    wb_stb_i,
    wb_we_i,
    write_enable_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rst_i;
 input wb_stb_i;
 input wb_we_i;
 input write_enable_i;
 input [5:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire \bit_sel[0] ;
 wire \bit_sel[10] ;
 wire \bit_sel[11] ;
 wire \bit_sel[12] ;
 wire \bit_sel[13] ;
 wire \bit_sel[14] ;
 wire \bit_sel[15] ;
 wire \bit_sel[16] ;
 wire \bit_sel[17] ;
 wire \bit_sel[18] ;
 wire \bit_sel[19] ;
 wire \bit_sel[1] ;
 wire \bit_sel[20] ;
 wire \bit_sel[21] ;
 wire \bit_sel[22] ;
 wire \bit_sel[23] ;
 wire \bit_sel[24] ;
 wire \bit_sel[25] ;
 wire \bit_sel[26] ;
 wire \bit_sel[27] ;
 wire \bit_sel[28] ;
 wire \bit_sel[29] ;
 wire \bit_sel[2] ;
 wire \bit_sel[30] ;
 wire \bit_sel[31] ;
 wire \bit_sel[32] ;
 wire \bit_sel[33] ;
 wire \bit_sel[34] ;
 wire \bit_sel[35] ;
 wire \bit_sel[36] ;
 wire \bit_sel[37] ;
 wire \bit_sel[38] ;
 wire \bit_sel[39] ;
 wire \bit_sel[3] ;
 wire \bit_sel[40] ;
 wire \bit_sel[41] ;
 wire \bit_sel[42] ;
 wire \bit_sel[43] ;
 wire \bit_sel[44] ;
 wire \bit_sel[45] ;
 wire \bit_sel[46] ;
 wire \bit_sel[47] ;
 wire \bit_sel[48] ;
 wire \bit_sel[49] ;
 wire \bit_sel[4] ;
 wire \bit_sel[50] ;
 wire \bit_sel[51] ;
 wire \bit_sel[52] ;
 wire \bit_sel[53] ;
 wire \bit_sel[54] ;
 wire \bit_sel[55] ;
 wire \bit_sel[56] ;
 wire \bit_sel[57] ;
 wire \bit_sel[58] ;
 wire \bit_sel[59] ;
 wire \bit_sel[5] ;
 wire \bit_sel[60] ;
 wire \bit_sel[61] ;
 wire \bit_sel[62] ;
 wire \bit_sel[63] ;
 wire \bit_sel[6] ;
 wire \bit_sel[7] ;
 wire \bit_sel[8] ;
 wire \bit_sel[9] ;
 wire \bit_sel_reg[0] ;
 wire \bit_sel_reg[10] ;
 wire \bit_sel_reg[11] ;
 wire \bit_sel_reg[12] ;
 wire \bit_sel_reg[13] ;
 wire \bit_sel_reg[14] ;
 wire \bit_sel_reg[15] ;
 wire \bit_sel_reg[16] ;
 wire \bit_sel_reg[17] ;
 wire \bit_sel_reg[18] ;
 wire \bit_sel_reg[19] ;
 wire \bit_sel_reg[1] ;
 wire \bit_sel_reg[20] ;
 wire \bit_sel_reg[21] ;
 wire \bit_sel_reg[22] ;
 wire \bit_sel_reg[23] ;
 wire \bit_sel_reg[24] ;
 wire \bit_sel_reg[25] ;
 wire \bit_sel_reg[26] ;
 wire \bit_sel_reg[27] ;
 wire \bit_sel_reg[28] ;
 wire \bit_sel_reg[29] ;
 wire \bit_sel_reg[2] ;
 wire \bit_sel_reg[30] ;
 wire \bit_sel_reg[31] ;
 wire \bit_sel_reg[32] ;
 wire \bit_sel_reg[33] ;
 wire \bit_sel_reg[34] ;
 wire \bit_sel_reg[35] ;
 wire \bit_sel_reg[36] ;
 wire \bit_sel_reg[37] ;
 wire \bit_sel_reg[38] ;
 wire \bit_sel_reg[39] ;
 wire \bit_sel_reg[3] ;
 wire \bit_sel_reg[40] ;
 wire \bit_sel_reg[41] ;
 wire \bit_sel_reg[42] ;
 wire \bit_sel_reg[43] ;
 wire \bit_sel_reg[44] ;
 wire \bit_sel_reg[45] ;
 wire \bit_sel_reg[46] ;
 wire \bit_sel_reg[47] ;
 wire \bit_sel_reg[48] ;
 wire \bit_sel_reg[49] ;
 wire \bit_sel_reg[4] ;
 wire \bit_sel_reg[50] ;
 wire \bit_sel_reg[51] ;
 wire \bit_sel_reg[52] ;
 wire \bit_sel_reg[53] ;
 wire \bit_sel_reg[54] ;
 wire \bit_sel_reg[55] ;
 wire \bit_sel_reg[56] ;
 wire \bit_sel_reg[57] ;
 wire \bit_sel_reg[58] ;
 wire \bit_sel_reg[59] ;
 wire \bit_sel_reg[5] ;
 wire \bit_sel_reg[60] ;
 wire \bit_sel_reg[61] ;
 wire \bit_sel_reg[62] ;
 wire \bit_sel_reg[63] ;
 wire \bit_sel_reg[6] ;
 wire \bit_sel_reg[7] ;
 wire \bit_sel_reg[8] ;
 wire \bit_sel_reg[9] ;
 wire \col_prog_n[0] ;
 wire \col_prog_n[10] ;
 wire \col_prog_n[11] ;
 wire \col_prog_n[12] ;
 wire \col_prog_n[13] ;
 wire \col_prog_n[14] ;
 wire \col_prog_n[15] ;
 wire \col_prog_n[16] ;
 wire \col_prog_n[17] ;
 wire \col_prog_n[18] ;
 wire \col_prog_n[19] ;
 wire \col_prog_n[1] ;
 wire \col_prog_n[20] ;
 wire \col_prog_n[21] ;
 wire \col_prog_n[22] ;
 wire \col_prog_n[23] ;
 wire \col_prog_n[24] ;
 wire \col_prog_n[25] ;
 wire \col_prog_n[26] ;
 wire \col_prog_n[27] ;
 wire \col_prog_n[28] ;
 wire \col_prog_n[29] ;
 wire \col_prog_n[2] ;
 wire \col_prog_n[30] ;
 wire \col_prog_n[31] ;
 wire \col_prog_n[3] ;
 wire \col_prog_n[4] ;
 wire \col_prog_n[5] ;
 wire \col_prog_n[6] ;
 wire \col_prog_n[7] ;
 wire \col_prog_n[8] ;
 wire \col_prog_n[9] ;
 wire \col_prog_n_reg[0] ;
 wire \col_prog_n_reg[10] ;
 wire \col_prog_n_reg[11] ;
 wire \col_prog_n_reg[12] ;
 wire \col_prog_n_reg[13] ;
 wire \col_prog_n_reg[14] ;
 wire \col_prog_n_reg[15] ;
 wire \col_prog_n_reg[16] ;
 wire \col_prog_n_reg[17] ;
 wire \col_prog_n_reg[18] ;
 wire \col_prog_n_reg[19] ;
 wire \col_prog_n_reg[1] ;
 wire \col_prog_n_reg[20] ;
 wire \col_prog_n_reg[21] ;
 wire \col_prog_n_reg[22] ;
 wire \col_prog_n_reg[23] ;
 wire \col_prog_n_reg[24] ;
 wire \col_prog_n_reg[25] ;
 wire \col_prog_n_reg[26] ;
 wire \col_prog_n_reg[27] ;
 wire \col_prog_n_reg[28] ;
 wire \col_prog_n_reg[29] ;
 wire \col_prog_n_reg[2] ;
 wire \col_prog_n_reg[30] ;
 wire \col_prog_n_reg[31] ;
 wire \col_prog_n_reg[3] ;
 wire \col_prog_n_reg[4] ;
 wire \col_prog_n_reg[5] ;
 wire \col_prog_n_reg[6] ;
 wire \col_prog_n_reg[7] ;
 wire \col_prog_n_reg[8] ;
 wire \col_prog_n_reg[9] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \efuse_out[0] ;
 wire \efuse_out[10] ;
 wire \efuse_out[11] ;
 wire \efuse_out[12] ;
 wire \efuse_out[13] ;
 wire \efuse_out[14] ;
 wire \efuse_out[15] ;
 wire \efuse_out[16] ;
 wire \efuse_out[17] ;
 wire \efuse_out[18] ;
 wire \efuse_out[19] ;
 wire \efuse_out[1] ;
 wire \efuse_out[20] ;
 wire \efuse_out[21] ;
 wire \efuse_out[22] ;
 wire \efuse_out[23] ;
 wire \efuse_out[24] ;
 wire \efuse_out[25] ;
 wire \efuse_out[26] ;
 wire \efuse_out[27] ;
 wire \efuse_out[28] ;
 wire \efuse_out[29] ;
 wire \efuse_out[2] ;
 wire \efuse_out[30] ;
 wire \efuse_out[31] ;
 wire \efuse_out[3] ;
 wire \efuse_out[4] ;
 wire \efuse_out[5] ;
 wire \efuse_out[6] ;
 wire \efuse_out[7] ;
 wire \efuse_out[8] ;
 wire \efuse_out[9] ;
 wire one;
 wire preset_n;
 wire preset_n_reg;
 wire sense;
 wire sense_del;
 wire sense_reg;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0524_ (.I(preset_n_reg),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0525_ (.I(\col_prog_n_reg[31] ),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0526_ (.I(\state[3] ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0527_ (.I(\col_prog_n_reg[30] ),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0528_ (.I(\col_prog_n_reg[29] ),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0529_ (.I(\col_prog_n_reg[28] ),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0530_ (.I(\col_prog_n_reg[27] ),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0531_ (.I(\col_prog_n_reg[26] ),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0532_ (.I(\col_prog_n_reg[25] ),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0533_ (.I(\col_prog_n_reg[24] ),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0534_ (.I(\col_prog_n_reg[23] ),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0535_ (.I(\col_prog_n_reg[22] ),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0536_ (.I(\col_prog_n_reg[21] ),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0537_ (.I(\col_prog_n_reg[20] ),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0538_ (.I(\col_prog_n_reg[19] ),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0539_ (.I(\col_prog_n_reg[18] ),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0540_ (.I(\col_prog_n_reg[17] ),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0541_ (.I(\col_prog_n_reg[16] ),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0542_ (.I(\col_prog_n_reg[15] ),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0543_ (.I(\col_prog_n_reg[14] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0544_ (.I(\col_prog_n_reg[13] ),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0545_ (.I(\col_prog_n_reg[12] ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0546_ (.I(\col_prog_n_reg[11] ),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0547_ (.I(\col_prog_n_reg[10] ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0548_ (.I(\col_prog_n_reg[9] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0549_ (.I(\col_prog_n_reg[8] ),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0550_ (.I(\col_prog_n_reg[7] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0551_ (.I(\col_prog_n_reg[6] ),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0552_ (.I(\col_prog_n_reg[5] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0553_ (.I(\col_prog_n_reg[4] ),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0554_ (.I(\col_prog_n_reg[3] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0555_ (.I(\col_prog_n_reg[2] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0556_ (.I(\col_prog_n_reg[1] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0557_ (.I(\col_prog_n_reg[0] ),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0558_ (.I(\counter[9] ),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0559_ (.I(\counter[8] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0560_ (.I(\counter[7] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0561_ (.I(\counter[6] ),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0562_ (.I(\counter[5] ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0563_ (.I(\counter[4] ),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0564_ (.I(\counter[3] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0565_ (.I(\counter[2] ),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0566_ (.I(\counter[1] ),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0567_ (.I(net47),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0568_ (.I(net90),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0569_ (.I(\state[0] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0570_ (.I(net6),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0571_ (.I(net2),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0572_ (.I(net1),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0573_ (.I(net4),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0574_ (.I(net5),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0575_ (.I(net92),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0576_ (.A1(net7),
    .A2(net45),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0577_ (.A1(net46),
    .A2(\state[0] ),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0578_ (.A1(net47),
    .A2(_0340_),
    .B(\state[0] ),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0579_ (.A1(net47),
    .A2(net46),
    .A3(_0340_),
    .B(\state[0] ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0580_ (.A1(\state[2] ),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0581_ (.A1(net47),
    .A2(net46),
    .A3(_0334_),
    .A4(_0340_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0582_ (.A1(_0289_),
    .A2(_0000_),
    .B(_0344_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0583_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0584_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .A4(\counter[0] ),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0585_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .A3(\counter[5] ),
    .A4(\counter[4] ),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0586_ (.A1(_0346_),
    .A2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0587_ (.A1(\counter[9] ),
    .A2(\counter[8] ),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0588_ (.A1(_0291_),
    .A2(_0346_),
    .A3(_0347_),
    .A4(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0589_ (.A1(\state[3] ),
    .A2(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0590_ (.A1(net44),
    .A2(net32),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0591_ (.A1(_0290_),
    .A2(net88),
    .B1(net84),
    .B2(_0352_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0592_ (.A1(net44),
    .A2(net31),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0593_ (.A1(net88),
    .A2(_0292_),
    .B1(net84),
    .B2(_0353_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0594_ (.A1(net44),
    .A2(net29),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0595_ (.A1(net88),
    .A2(_0293_),
    .B1(net84),
    .B2(_0354_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0596_ (.A1(net44),
    .A2(net28),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0597_ (.A1(net88),
    .A2(_0294_),
    .B1(net84),
    .B2(_0355_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0598_ (.A1(net44),
    .A2(net27),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0599_ (.A1(net88),
    .A2(_0295_),
    .B1(net84),
    .B2(_0356_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0600_ (.A1(net44),
    .A2(net26),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0601_ (.A1(_0291_),
    .A2(_0296_),
    .B1(net84),
    .B2(_0357_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0602_ (.A1(net44),
    .A2(net25),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0603_ (.A1(_0291_),
    .A2(_0297_),
    .B1(_0351_),
    .B2(_0358_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0604_ (.A1(net44),
    .A2(net24),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0605_ (.A1(_0291_),
    .A2(_0298_),
    .B1(_0351_),
    .B2(_0359_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0606_ (.A1(net43),
    .A2(net23),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0607_ (.A1(_0291_),
    .A2(_0299_),
    .B1(_0351_),
    .B2(_0360_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0608_ (.A1(net43),
    .A2(net22),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0609_ (.A1(_0291_),
    .A2(_0300_),
    .B1(_0351_),
    .B2(_0361_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0610_ (.A1(net43),
    .A2(net21),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0611_ (.A1(_0291_),
    .A2(_0301_),
    .B1(_0351_),
    .B2(_0362_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0612_ (.A1(net43),
    .A2(net20),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0613_ (.A1(_0291_),
    .A2(_0302_),
    .B1(_0351_),
    .B2(_0363_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0614_ (.A1(net43),
    .A2(net18),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0615_ (.A1(_0291_),
    .A2(_0303_),
    .B1(_0351_),
    .B2(_0364_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0616_ (.A1(net43),
    .A2(net17),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0617_ (.A1(_0291_),
    .A2(_0304_),
    .B1(_0351_),
    .B2(_0365_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0618_ (.A1(net43),
    .A2(net16),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0619_ (.A1(_0291_),
    .A2(_0305_),
    .B1(_0351_),
    .B2(_0366_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0620_ (.A1(net43),
    .A2(net15),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0621_ (.A1(net88),
    .A2(_0306_),
    .B1(net84),
    .B2(_0367_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0622_ (.A1(net42),
    .A2(net14),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0623_ (.A1(_0291_),
    .A2(_0307_),
    .B1(_0351_),
    .B2(_0368_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0624_ (.A1(net42),
    .A2(net13),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0625_ (.A1(net88),
    .A2(_0308_),
    .B1(net84),
    .B2(_0369_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0626_ (.A1(net42),
    .A2(net12),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0627_ (.A1(net88),
    .A2(_0309_),
    .B1(net84),
    .B2(_0370_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0628_ (.A1(net42),
    .A2(net11),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0629_ (.A1(net88),
    .A2(_0310_),
    .B1(net84),
    .B2(_0371_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0630_ (.A1(net42),
    .A2(net10),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0631_ (.A1(net88),
    .A2(_0311_),
    .B1(net84),
    .B2(_0372_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0632_ (.A1(net42),
    .A2(net9),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0633_ (.A1(net88),
    .A2(_0312_),
    .B1(net84),
    .B2(_0373_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0634_ (.A1(net42),
    .A2(net39),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0635_ (.A1(_0291_),
    .A2(_0313_),
    .B1(_0351_),
    .B2(_0374_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0636_ (.A1(net42),
    .A2(net38),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0637_ (.A1(net88),
    .A2(_0314_),
    .B1(net84),
    .B2(_0375_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0638_ (.A1(net41),
    .A2(net37),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0639_ (.A1(net88),
    .A2(_0315_),
    .B1(net84),
    .B2(_0376_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0640_ (.A1(net41),
    .A2(net36),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0641_ (.A1(net88),
    .A2(_0316_),
    .B1(net84),
    .B2(_0377_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0642_ (.A1(net41),
    .A2(net35),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0643_ (.A1(net88),
    .A2(_0317_),
    .B1(net84),
    .B2(_0378_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0644_ (.A1(net41),
    .A2(net34),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0645_ (.A1(net88),
    .A2(_0318_),
    .B1(net84),
    .B2(_0379_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0646_ (.A1(net41),
    .A2(net33),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0647_ (.A1(net88),
    .A2(_0319_),
    .B1(net84),
    .B2(_0380_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0648_ (.A1(net41),
    .A2(net30),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0649_ (.A1(net88),
    .A2(_0320_),
    .B1(net84),
    .B2(_0381_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0650_ (.A1(net41),
    .A2(net19),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0651_ (.A1(net88),
    .A2(_0321_),
    .B1(net84),
    .B2(_0382_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0652_ (.A1(net41),
    .A2(net8),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0653_ (.A1(net88),
    .A2(_0322_),
    .B1(net84),
    .B2(_0383_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0654_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0655_ (.A1(\bit_sel_reg[63] ),
    .A2(net86),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0656_ (.A1(net2),
    .A2(net1),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0657_ (.A1(net2),
    .A2(net1),
    .A3(net3),
    .A4(net4),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0658_ (.A1(net5),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0659_ (.A1(net47),
    .A2(_0340_),
    .A3(_0341_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0660_ (.A1(net47),
    .A2(_0340_),
    .A3(_0341_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0661_ (.A1(\state[2] ),
    .A2(_0389_),
    .B(net6),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0662_ (.A1(_0388_),
    .A2(net82),
    .B(_0385_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0663_ (.A1(\bit_sel_reg[62] ),
    .A2(_0384_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0664_ (.A1(_0336_),
    .A2(net1),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0665_ (.A1(net3),
    .A2(net4),
    .A3(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0666_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0393_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0667_ (.A1(_0391_),
    .A2(_0395_),
    .B(_0392_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0668_ (.A1(\bit_sel_reg[61] ),
    .A2(_0384_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0669_ (.A1(net2),
    .A2(_0337_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0670_ (.A1(net3),
    .A2(net4),
    .A3(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0671_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0397_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0672_ (.A1(_0391_),
    .A2(_0399_),
    .B(_0396_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0673_ (.A1(\bit_sel_reg[60] ),
    .A2(net86),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0674_ (.A1(net2),
    .A2(net1),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0675_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0676_ (.A1(net83),
    .A2(_0402_),
    .B(_0400_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0677_ (.A1(\bit_sel_reg[59] ),
    .A2(net86),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0678_ (.A1(net3),
    .A2(_0386_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0679_ (.A1(net4),
    .A2(net5),
    .A3(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0680_ (.A1(net83),
    .A2(_0405_),
    .B(_0403_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0681_ (.A1(\bit_sel_reg[58] ),
    .A2(net87),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0682_ (.A1(_0336_),
    .A2(net1),
    .A3(net3),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0683_ (.A1(net4),
    .A2(net5),
    .A3(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0684_ (.A1(net83),
    .A2(_0408_),
    .B(_0406_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0685_ (.A1(\bit_sel_reg[57] ),
    .A2(net87),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0686_ (.A1(net2),
    .A2(_0337_),
    .A3(net3),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0687_ (.A1(net4),
    .A2(net5),
    .A3(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0688_ (.A1(_0391_),
    .A2(_0411_),
    .B(_0409_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0689_ (.A1(\bit_sel_reg[56] ),
    .A2(net86),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0690_ (.A1(net2),
    .A2(net1),
    .A3(net3),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0691_ (.A1(net4),
    .A2(net5),
    .A3(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0692_ (.A1(net83),
    .A2(_0414_),
    .B(_0412_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0693_ (.A1(\bit_sel_reg[55] ),
    .A2(net87),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0694_ (.A1(net2),
    .A2(net1),
    .A3(net3),
    .A4(_0338_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0695_ (.A1(net5),
    .A2(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0696_ (.A1(net82),
    .A2(_0417_),
    .B(_0415_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0697_ (.A1(\bit_sel_reg[54] ),
    .A2(_0384_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0698_ (.A1(net3),
    .A2(_0338_),
    .A3(net5),
    .A4(_0393_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0699_ (.A1(_0391_),
    .A2(_0419_),
    .B(_0418_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0700_ (.A1(\bit_sel_reg[53] ),
    .A2(_0384_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0701_ (.A1(net3),
    .A2(_0338_),
    .A3(net5),
    .A4(_0397_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0702_ (.A1(_0391_),
    .A2(_0421_),
    .B(_0420_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0703_ (.A1(\bit_sel_reg[52] ),
    .A2(net86),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0704_ (.A1(net3),
    .A2(_0338_),
    .A3(net5),
    .A4(_0401_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0705_ (.A1(net83),
    .A2(_0423_),
    .B(_0422_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0706_ (.A1(\bit_sel_reg[51] ),
    .A2(net87),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0707_ (.A1(net3),
    .A2(net4),
    .A3(_0386_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0708_ (.A1(net5),
    .A2(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0709_ (.A1(net82),
    .A2(_0426_),
    .B(_0424_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0710_ (.A1(\bit_sel_reg[50] ),
    .A2(net86),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0711_ (.A1(_0336_),
    .A2(net1),
    .A3(net3),
    .A4(net4),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0712_ (.A1(net5),
    .A2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0713_ (.A1(net82),
    .A2(_0429_),
    .B(_0427_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0714_ (.A1(\bit_sel_reg[49] ),
    .A2(net86),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0715_ (.A1(net2),
    .A2(_0337_),
    .A3(net3),
    .A4(net4),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0716_ (.A1(net5),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0717_ (.A1(net83),
    .A2(_0432_),
    .B(_0430_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0718_ (.A1(\bit_sel_reg[48] ),
    .A2(net86),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0719_ (.A1(_0338_),
    .A2(_0413_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0720_ (.A1(net5),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0721_ (.A1(net82),
    .A2(_0435_),
    .B(_0433_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0722_ (.A1(\bit_sel_reg[47] ),
    .A2(net86),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0723_ (.A1(_0339_),
    .A2(_0387_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0724_ (.A1(net83),
    .A2(_0437_),
    .B(_0436_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0725_ (.A1(\bit_sel_reg[46] ),
    .A2(_0384_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0726_ (.A1(net5),
    .A2(_0391_),
    .A3(_0394_),
    .B(_0438_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0727_ (.A1(\bit_sel_reg[45] ),
    .A2(_0384_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0728_ (.A1(net5),
    .A2(_0391_),
    .A3(_0398_),
    .B(_0439_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0729_ (.A1(\bit_sel_reg[44] ),
    .A2(net87),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0730_ (.A1(net3),
    .A2(net4),
    .A3(_0339_),
    .A4(_0401_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0731_ (.A1(net82),
    .A2(_0441_),
    .B(_0440_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0732_ (.A1(\bit_sel_reg[43] ),
    .A2(net87),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0733_ (.A1(net4),
    .A2(_0339_),
    .A3(_0404_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0734_ (.A1(net82),
    .A2(_0443_),
    .B(_0442_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0735_ (.A1(\bit_sel_reg[42] ),
    .A2(net87),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0736_ (.A1(net4),
    .A2(_0339_),
    .A3(_0407_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0737_ (.A1(_0391_),
    .A2(_0445_),
    .B(_0444_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0738_ (.A1(\bit_sel_reg[41] ),
    .A2(net87),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0739_ (.A1(net4),
    .A2(_0339_),
    .A3(_0410_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0740_ (.A1(net83),
    .A2(_0447_),
    .B(_0446_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0741_ (.A1(\bit_sel_reg[40] ),
    .A2(net87),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0742_ (.A1(net4),
    .A2(_0339_),
    .A3(_0413_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0743_ (.A1(net82),
    .A2(_0449_),
    .B(_0448_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0744_ (.A1(\bit_sel_reg[39] ),
    .A2(net87),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0745_ (.A1(_0339_),
    .A2(_0416_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0746_ (.A1(net82),
    .A2(_0451_),
    .B(_0450_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0747_ (.A1(\bit_sel_reg[38] ),
    .A2(net87),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0748_ (.A1(net3),
    .A2(_0338_),
    .A3(_0339_),
    .A4(_0393_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0749_ (.A1(net83),
    .A2(_0453_),
    .B(_0452_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0750_ (.A1(\bit_sel_reg[37] ),
    .A2(_0384_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0751_ (.A1(net3),
    .A2(_0338_),
    .A3(_0339_),
    .A4(_0397_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0752_ (.A1(_0391_),
    .A2(_0455_),
    .B(_0454_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0753_ (.A1(\bit_sel_reg[36] ),
    .A2(net86),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0754_ (.A1(net3),
    .A2(_0338_),
    .A3(_0339_),
    .A4(_0401_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0755_ (.A1(net83),
    .A2(_0457_),
    .B(_0456_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0756_ (.A1(\bit_sel_reg[35] ),
    .A2(net87),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0757_ (.A1(_0339_),
    .A2(_0425_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0758_ (.A1(net82),
    .A2(_0459_),
    .B(_0458_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0759_ (.A1(\bit_sel_reg[34] ),
    .A2(net86),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0760_ (.A1(_0339_),
    .A2(_0428_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0761_ (.A1(net83),
    .A2(_0461_),
    .B(_0460_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0762_ (.A1(\bit_sel_reg[33] ),
    .A2(net87),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0763_ (.A1(_0339_),
    .A2(_0431_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0764_ (.A1(net82),
    .A2(_0463_),
    .B(_0462_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0765_ (.A1(\bit_sel_reg[32] ),
    .A2(net87),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0766_ (.A1(_0339_),
    .A2(_0434_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0767_ (.A1(net82),
    .A2(_0465_),
    .B(_0464_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0768_ (.A1(\bit_sel_reg[31] ),
    .A2(net86),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0769_ (.A1(\state[2] ),
    .A2(_0389_),
    .B(_0335_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0770_ (.A1(_0388_),
    .A2(net80),
    .B(_0466_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0771_ (.A1(\bit_sel_reg[30] ),
    .A2(_0384_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0772_ (.A1(_0395_),
    .A2(_0467_),
    .B(_0468_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0773_ (.A1(\bit_sel_reg[29] ),
    .A2(_0384_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0774_ (.A1(_0399_),
    .A2(_0467_),
    .B(_0469_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0775_ (.A1(\bit_sel_reg[28] ),
    .A2(net86),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0776_ (.A1(_0402_),
    .A2(net81),
    .B(_0470_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0777_ (.A1(\bit_sel_reg[27] ),
    .A2(net86),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0778_ (.A1(_0405_),
    .A2(net80),
    .B(_0471_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0779_ (.A1(\bit_sel_reg[26] ),
    .A2(net87),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0780_ (.A1(_0408_),
    .A2(_0467_),
    .B(_0472_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0781_ (.A1(\bit_sel_reg[25] ),
    .A2(net87),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0782_ (.A1(_0411_),
    .A2(net81),
    .B(_0473_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0783_ (.A1(\bit_sel_reg[24] ),
    .A2(net86),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0784_ (.A1(_0414_),
    .A2(net80),
    .B(_0474_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0785_ (.A1(\bit_sel_reg[23] ),
    .A2(net87),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0786_ (.A1(_0417_),
    .A2(net80),
    .B(_0475_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0787_ (.A1(\bit_sel_reg[22] ),
    .A2(_0384_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0788_ (.A1(_0419_),
    .A2(net81),
    .B(_0476_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0789_ (.A1(\bit_sel_reg[21] ),
    .A2(_0384_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0790_ (.A1(_0421_),
    .A2(net81),
    .B(_0477_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0791_ (.A1(\bit_sel_reg[20] ),
    .A2(net86),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0792_ (.A1(_0423_),
    .A2(net81),
    .B(_0478_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0793_ (.A1(\bit_sel_reg[19] ),
    .A2(net87),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0794_ (.A1(_0426_),
    .A2(net80),
    .B(_0479_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0795_ (.A1(\bit_sel_reg[18] ),
    .A2(net86),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0796_ (.A1(_0429_),
    .A2(net80),
    .B(_0480_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0797_ (.A1(\bit_sel_reg[17] ),
    .A2(net86),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0798_ (.A1(_0432_),
    .A2(net81),
    .B(_0481_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0799_ (.A1(\bit_sel_reg[16] ),
    .A2(net86),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0800_ (.A1(_0435_),
    .A2(net80),
    .B(_0482_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0801_ (.A1(\bit_sel_reg[15] ),
    .A2(net86),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0802_ (.A1(_0437_),
    .A2(net80),
    .B(_0483_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0803_ (.A1(\bit_sel_reg[14] ),
    .A2(_0384_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0804_ (.A1(net5),
    .A2(_0394_),
    .A3(_0467_),
    .B(_0484_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0805_ (.A1(\bit_sel_reg[13] ),
    .A2(_0384_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0806_ (.A1(net5),
    .A2(_0398_),
    .A3(_0467_),
    .B(_0485_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0807_ (.A1(\bit_sel_reg[12] ),
    .A2(net87),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0808_ (.A1(_0441_),
    .A2(net81),
    .B(_0486_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0809_ (.A1(\bit_sel_reg[11] ),
    .A2(net87),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0810_ (.A1(_0443_),
    .A2(net81),
    .B(_0487_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0811_ (.A1(\bit_sel_reg[10] ),
    .A2(net87),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0812_ (.A1(_0445_),
    .A2(_0467_),
    .B(_0488_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0813_ (.A1(\bit_sel_reg[9] ),
    .A2(net87),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0814_ (.A1(_0447_),
    .A2(_0467_),
    .B(_0489_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0815_ (.A1(\bit_sel_reg[8] ),
    .A2(net87),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0816_ (.A1(_0449_),
    .A2(net81),
    .B(_0490_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0817_ (.A1(\bit_sel_reg[7] ),
    .A2(net87),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0818_ (.A1(_0451_),
    .A2(net80),
    .B(_0491_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0819_ (.A1(\bit_sel_reg[6] ),
    .A2(net87),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0820_ (.A1(_0453_),
    .A2(_0467_),
    .B(_0492_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0821_ (.A1(\bit_sel_reg[5] ),
    .A2(_0384_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0822_ (.A1(_0455_),
    .A2(net81),
    .B(_0493_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0823_ (.A1(\bit_sel_reg[4] ),
    .A2(net86),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0824_ (.A1(_0457_),
    .A2(net81),
    .B(_0494_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0825_ (.A1(\bit_sel_reg[3] ),
    .A2(net87),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0826_ (.A1(_0459_),
    .A2(net80),
    .B(_0495_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0827_ (.A1(\bit_sel_reg[2] ),
    .A2(net86),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0828_ (.A1(_0461_),
    .A2(net80),
    .B(_0496_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0829_ (.A1(\bit_sel_reg[1] ),
    .A2(net87),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0830_ (.A1(_0463_),
    .A2(net80),
    .B(_0497_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0831_ (.A1(\bit_sel_reg[0] ),
    .A2(net87),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0832_ (.A1(_0465_),
    .A2(net80),
    .B(_0498_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0833_ (.A1(net47),
    .A2(_0340_),
    .A3(_0341_),
    .B1(\state[0] ),
    .B2(_0291_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0834_ (.A1(_0350_),
    .A2(net85),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0835_ (.A1(_0350_),
    .A2(net85),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0836_ (.A1(_0324_),
    .A2(_0348_),
    .A3(_0350_),
    .A4(_0499_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0837_ (.A1(\state[3] ),
    .A2(_0390_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0838_ (.A1(\state[3] ),
    .A2(_0390_),
    .B1(_0502_),
    .B2(_0323_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0839_ (.A1(_0348_),
    .A2(_0499_),
    .B(_0324_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0840_ (.A1(_0502_),
    .A2(_0503_),
    .A3(_0504_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0841_ (.A1(\counter[4] ),
    .A2(_0346_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0842_ (.A1(\counter[5] ),
    .A2(\counter[4] ),
    .A3(_0346_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0843_ (.A1(\counter[6] ),
    .A2(\counter[5] ),
    .A3(\counter[4] ),
    .A4(_0346_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0844_ (.A1(_0291_),
    .A2(_0507_),
    .B(net85),
    .C(_0350_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0845_ (.A1(\state[3] ),
    .A2(_0350_),
    .A3(net85),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0846_ (.A1(\state[3] ),
    .A2(_0350_),
    .A3(net85),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0847_ (.A1(\counter[7] ),
    .A2(_0507_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0848_ (.A1(_0325_),
    .A2(_0508_),
    .B1(_0509_),
    .B2(_0511_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0849_ (.A1(_0350_),
    .A2(net85),
    .A3(_0506_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0850_ (.A1(_0326_),
    .A2(_0512_),
    .B(_0508_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0851_ (.A1(_0350_),
    .A2(net85),
    .A3(_0505_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0852_ (.A1(_0291_),
    .A2(_0506_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0853_ (.A1(_0327_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0501_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0854_ (.A1(\state[3] ),
    .A2(_0346_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0855_ (.A1(_0350_),
    .A2(net85),
    .A3(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0856_ (.A1(_0350_),
    .A2(net85),
    .A3(_0515_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0857_ (.A1(\state[3] ),
    .A2(_0350_),
    .A3(net85),
    .A4(_0505_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0858_ (.A1(_0328_),
    .A2(_0516_),
    .B(_0518_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0859_ (.A1(_0330_),
    .A2(_0345_),
    .A3(_0350_),
    .A4(net85),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0860_ (.A1(_0329_),
    .A2(_0519_),
    .B(_0517_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0861_ (.A1(_0330_),
    .A2(_0345_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0862_ (.A1(_0330_),
    .A2(_0500_),
    .B1(_0510_),
    .B2(_0520_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0863_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0864_ (.A1(_0331_),
    .A2(_0500_),
    .B1(_0510_),
    .B2(_0521_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0865_ (.I0(_0509_),
    .I1(_0501_),
    .S(\counter[0] ),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0866_ (.A1(_0333_),
    .A2(_0334_),
    .B1(_0350_),
    .B2(\state[3] ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0867_ (.A1(\state[3] ),
    .A2(_0333_),
    .B1(_0522_),
    .B2(_0332_),
    .C(_0350_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0868_ (.I0(net72),
    .I1(\efuse_out[31] ),
    .S(net89),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0869_ (.I0(net71),
    .I1(\efuse_out[30] ),
    .S(net89),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0870_ (.I0(net69),
    .I1(\efuse_out[29] ),
    .S(net89),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0871_ (.I0(net68),
    .I1(\efuse_out[28] ),
    .S(net90),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0872_ (.I0(net67),
    .I1(\efuse_out[27] ),
    .S(net90),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0873_ (.I0(net66),
    .I1(\efuse_out[26] ),
    .S(net90),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0874_ (.I0(net65),
    .I1(\efuse_out[25] ),
    .S(net90),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0875_ (.I0(net64),
    .I1(\efuse_out[24] ),
    .S(net90),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0876_ (.I0(net63),
    .I1(\efuse_out[23] ),
    .S(\state[1] ),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0877_ (.I0(net62),
    .I1(\efuse_out[22] ),
    .S(\state[1] ),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0878_ (.I0(net61),
    .I1(\efuse_out[21] ),
    .S(\state[1] ),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0879_ (.I0(net60),
    .I1(\efuse_out[20] ),
    .S(net89),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0880_ (.I0(net58),
    .I1(\efuse_out[19] ),
    .S(net90),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0881_ (.I0(net57),
    .I1(\efuse_out[18] ),
    .S(net89),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0882_ (.I0(net56),
    .I1(\efuse_out[17] ),
    .S(net89),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0883_ (.I0(net55),
    .I1(\efuse_out[16] ),
    .S(net89),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0884_ (.I0(net54),
    .I1(\efuse_out[15] ),
    .S(net90),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0885_ (.I0(net53),
    .I1(\efuse_out[14] ),
    .S(net90),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0886_ (.I0(net52),
    .I1(\efuse_out[13] ),
    .S(net90),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0887_ (.I0(net51),
    .I1(\efuse_out[12] ),
    .S(net90),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0888_ (.I0(net50),
    .I1(\efuse_out[11] ),
    .S(net89),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0889_ (.I0(net49),
    .I1(\efuse_out[10] ),
    .S(net89),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0890_ (.I0(net79),
    .I1(\efuse_out[9] ),
    .S(net89),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0891_ (.I0(net78),
    .I1(\efuse_out[8] ),
    .S(net90),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0892_ (.I0(net77),
    .I1(\efuse_out[7] ),
    .S(net89),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0893_ (.I0(net76),
    .I1(\efuse_out[6] ),
    .S(net89),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0894_ (.I0(net75),
    .I1(\efuse_out[5] ),
    .S(\state[1] ),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0895_ (.I0(net74),
    .I1(\efuse_out[4] ),
    .S(net90),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0896_ (.I0(net73),
    .I1(\efuse_out[3] ),
    .S(net90),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0897_ (.I0(net70),
    .I1(\efuse_out[2] ),
    .S(net89),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0898_ (.I0(net59),
    .I1(\efuse_out[1] ),
    .S(net89),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0899_ (.I0(net48),
    .I1(\efuse_out[0] ),
    .S(net89),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0900_ (.A1(sense_reg),
    .A2(_0000_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0901_ (.A1(\state[1] ),
    .A2(_0343_),
    .B(_0523_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0902_ (.A1(_0351_),
    .A2(_0389_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0903_ (.A1(_0333_),
    .A2(_0342_),
    .A3(_0350_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0904_ (.I(net92),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0905_ (.I(net92),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0906_ (.I(net92),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0907_ (.I(net92),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0908_ (.I(net40),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0909_ (.I(net40),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0910_ (.I(net40),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0911_ (.I(net92),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0912_ (.I(net92),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0913_ (.I(net92),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0914_ (.I(net40),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0915_ (.I(net92),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0916_ (.I(net92),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0917_ (.I(net40),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0918_ (.I(net40),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0919_ (.I(net40),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0920_ (.I(net92),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0921_ (.I(net92),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0922_ (.I(net92),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0923_ (.I(net92),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0924_ (.I(net40),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0925_ (.I(net92),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0926_ (.I(net40),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0927_ (.I(net92),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0928_ (.I(net40),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0929_ (.I(net92),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0930_ (.I(net92),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0931_ (.I(net92),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0932_ (.I(net92),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0933_ (.I(net92),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0934_ (.I(net92),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0935_ (.I(net40),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0936_ (.I(net40),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0937_ (.I(net40),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0938_ (.I(net40),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0939_ (.I(net40),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0940_ (.I(net92),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0941_ (.I(net92),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0942_ (.I(net92),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0943_ (.I(net92),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0944_ (.I(net92),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0945_ (.I(net92),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0946_ (.I(net92),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0947_ (.I(net92),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0948_ (.I(net92),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0949_ (.I(net92),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0950_ (.I(net92),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0951_ (.I(net91),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0952_ (.I(net91),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0953_ (.I(net91),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0954_ (.I(net91),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0955_ (.I(net91),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0956_ (.I(net91),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0957_ (.I(net91),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0958_ (.I(net91),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0959_ (.I(net91),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0960_ (.I(net91),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0961_ (.I(net91),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0962_ (.I(net91),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0963_ (.I(net91),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0964_ (.I(net91),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0965_ (.I(net92),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0966_ (.I(net91),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0967_ (.I(net91),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0968_ (.I(net91),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0969_ (.I(net91),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0970_ (.I(net91),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0971_ (.I(net91),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0972_ (.I(net91),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0973_ (.I(net91),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0974_ (.I(net91),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0975_ (.I(net91),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0976_ (.I(net91),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0977_ (.I(net91),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0978_ (.I(net91),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0979_ (.I(net91),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0980_ (.I(net91),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0981_ (.I(net91),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0982_ (.I(net91),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0983_ (.I(net91),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0984_ (.I(net91),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0985_ (.I(net91),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0986_ (.I(net91),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0987_ (.I(net91),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0988_ (.I(net91),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0989_ (.I(net91),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0990_ (.I(net91),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0991_ (.I(net91),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0992_ (.I(net91),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0993_ (.I(net91),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0994_ (.I(net91),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0995_ (.I(net91),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0996_ (.I(net91),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0997_ (.I(net92),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0998_ (.I(net91),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0999_ (.I(net91),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1000_ (.I(net91),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1001_ (.I(net91),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1002_ (.I(net91),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1003_ (.I(net91),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1004_ (.I(net91),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1005_ (.I(net91),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1006_ (.I(net91),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1007_ (.I(net91),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1008_ (.I(net91),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1009_ (.I(net91),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1010_ (.I(net91),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1011_ (.I(net91),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1012_ (.I(net91),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1013_ (.I(net92),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1014_ (.I(net91),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1015_ (.I(net40),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1016_ (.I(net40),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1017_ (.I(net40),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1018_ (.I(net40),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1019_ (.I(net40),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1020_ (.I(net40),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1021_ (.I(net40),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1022_ (.I(net40),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1023_ (.I(net40),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1024_ (.I(net92),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1025_ (.I(net40),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1026_ (.I(net40),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1027_ (.I(net40),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1028_ (.I(net40),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1029_ (.I(net92),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1030_ (.I(net92),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1031_ (.I(net92),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1032_ (.I(net92),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1033_ (.I(net92),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1034_ (.I(net92),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1035_ (.I(net92),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1036_ (.I(net92),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1037_ (.I(net92),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1038_ (.I(net92),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1039_ (.I(net92),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1040_ (.I(net92),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1041_ (.I(net92),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1042_ (.I(net40),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1043_ (.I(net40),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1044_ (.I(net40),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1045_ (.I(net40),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1046_ (.I(net40),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1047_ (.I(net92),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1048_ (.D(_0001_),
    .SETN(_0003_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1049_ (.D(\state[2] ),
    .RN(_0004_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1050_ (.D(_0000_),
    .RN(_0005_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1051_ (.D(_0002_),
    .RN(_0006_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1052_ (.D(_0148_),
    .RN(_0007_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(sense_reg));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1053_ (.D(_0149_),
    .RN(_0008_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1054_ (.D(_0150_),
    .RN(_0009_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1055_ (.D(_0151_),
    .RN(_0010_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1056_ (.D(_0152_),
    .RN(_0011_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1057_ (.D(_0153_),
    .RN(_0012_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1058_ (.D(_0154_),
    .RN(_0013_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1059_ (.D(_0155_),
    .RN(_0014_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net76));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1060_ (.D(_0156_),
    .RN(_0015_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1061_ (.D(_0157_),
    .RN(_0016_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1062_ (.D(_0158_),
    .RN(_0017_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1063_ (.D(_0159_),
    .RN(_0018_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1064_ (.D(_0160_),
    .RN(_0019_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1065_ (.D(_0161_),
    .RN(_0020_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1066_ (.D(_0162_),
    .RN(_0021_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1067_ (.D(_0163_),
    .RN(_0022_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1068_ (.D(_0164_),
    .RN(_0023_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1069_ (.D(_0165_),
    .RN(_0024_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1070_ (.D(_0166_),
    .RN(_0025_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1071_ (.D(_0167_),
    .RN(_0026_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1072_ (.D(_0168_),
    .RN(_0027_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1073_ (.D(_0169_),
    .RN(_0028_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1074_ (.D(_0170_),
    .RN(_0029_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1075_ (.D(_0171_),
    .RN(_0030_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1076_ (.D(_0172_),
    .RN(_0031_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1077_ (.D(_0173_),
    .RN(_0032_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1078_ (.D(_0174_),
    .RN(_0033_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1079_ (.D(_0175_),
    .RN(_0034_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1080_ (.D(_0176_),
    .RN(_0035_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1081_ (.D(_0177_),
    .RN(_0036_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1082_ (.D(_0178_),
    .RN(_0037_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1083_ (.D(_0179_),
    .RN(_0038_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1084_ (.D(_0180_),
    .RN(_0039_),
    .CLK(clknet_4_1__leaf_wb_clk_i),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1085_ (.D(_0181_),
    .RN(_0040_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1086_ (.D(_0182_),
    .RN(_0041_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1087_ (.D(_0183_),
    .RN(_0042_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1088_ (.D(_0184_),
    .RN(_0043_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1089_ (.D(_0185_),
    .RN(_0044_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1090_ (.D(_0186_),
    .RN(_0045_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1091_ (.D(_0187_),
    .RN(_0046_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1092_ (.D(_0188_),
    .RN(_0047_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1093_ (.D(_0189_),
    .RN(_0048_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1094_ (.D(_0190_),
    .RN(_0049_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1095_ (.D(_0191_),
    .RN(_0050_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1096_ (.D(_0192_),
    .RN(_0051_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1097_ (.D(_0193_),
    .RN(_0052_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1098_ (.D(_0194_),
    .RN(_0053_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1099_ (.D(_0195_),
    .RN(_0054_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1100_ (.D(_0196_),
    .RN(_0055_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1101_ (.D(_0197_),
    .RN(_0056_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1102_ (.D(_0198_),
    .RN(_0057_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1103_ (.D(_0199_),
    .RN(_0058_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1104_ (.D(_0200_),
    .RN(_0059_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1105_ (.D(_0201_),
    .RN(_0060_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1106_ (.D(_0202_),
    .RN(_0061_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1107_ (.D(_0203_),
    .RN(_0062_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1108_ (.D(_0204_),
    .RN(_0063_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1109_ (.D(_0205_),
    .RN(_0064_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1110_ (.D(_0206_),
    .RN(_0065_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\bit_sel_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1111_ (.D(_0207_),
    .RN(_0066_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1112_ (.D(_0208_),
    .RN(_0067_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1113_ (.D(_0209_),
    .RN(_0068_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1114_ (.D(_0210_),
    .RN(_0069_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1115_ (.D(_0211_),
    .RN(_0070_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1116_ (.D(_0212_),
    .RN(_0071_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1117_ (.D(_0213_),
    .RN(_0072_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1118_ (.D(_0214_),
    .RN(_0073_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1119_ (.D(_0215_),
    .RN(_0074_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1120_ (.D(_0216_),
    .RN(_0075_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1121_ (.D(_0217_),
    .RN(_0076_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1122_ (.D(_0218_),
    .RN(_0077_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1123_ (.D(_0219_),
    .RN(_0078_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1124_ (.D(_0220_),
    .RN(_0079_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1125_ (.D(_0221_),
    .RN(_0080_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\bit_sel_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1126_ (.D(_0222_),
    .RN(_0081_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\bit_sel_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1127_ (.D(_0223_),
    .RN(_0082_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1128_ (.D(_0224_),
    .RN(_0083_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1129_ (.D(_0225_),
    .RN(_0084_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1130_ (.D(_0226_),
    .RN(_0085_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1131_ (.D(_0227_),
    .RN(_0086_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1132_ (.D(_0228_),
    .RN(_0087_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1133_ (.D(_0229_),
    .RN(_0088_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\bit_sel_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1134_ (.D(_0230_),
    .RN(_0089_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1135_ (.D(_0231_),
    .RN(_0090_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1136_ (.D(_0232_),
    .RN(_0091_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1137_ (.D(_0233_),
    .RN(_0092_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1138_ (.D(_0234_),
    .RN(_0093_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1139_ (.D(_0235_),
    .RN(_0094_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1140_ (.D(_0236_),
    .RN(_0095_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1141_ (.D(_0237_),
    .RN(_0096_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1142_ (.D(_0238_),
    .RN(_0097_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\bit_sel_reg[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1143_ (.D(_0239_),
    .RN(_0098_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1144_ (.D(_0240_),
    .RN(_0099_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1145_ (.D(_0241_),
    .RN(_0100_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1146_ (.D(_0242_),
    .RN(_0101_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1147_ (.D(_0243_),
    .RN(_0102_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1148_ (.D(_0244_),
    .RN(_0103_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1149_ (.D(_0245_),
    .RN(_0104_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1150_ (.D(_0246_),
    .RN(_0105_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\bit_sel_reg[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1151_ (.D(_0247_),
    .RN(_0106_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1152_ (.D(_0248_),
    .RN(_0107_),
    .CLK(clknet_4_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1153_ (.D(_0249_),
    .RN(_0108_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1154_ (.D(_0250_),
    .RN(_0109_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1155_ (.D(_0251_),
    .RN(_0110_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1156_ (.D(_0252_),
    .RN(_0111_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1157_ (.D(_0253_),
    .RN(_0112_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\bit_sel_reg[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1158_ (.D(_0254_),
    .RN(_0113_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\bit_sel_reg[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1159_ (.D(_0255_),
    .RN(_0114_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1160_ (.D(_0256_),
    .SETN(_0115_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1161_ (.D(_0257_),
    .SETN(_0116_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1162_ (.D(_0258_),
    .SETN(_0117_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1163_ (.D(_0259_),
    .SETN(_0118_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1164_ (.D(_0260_),
    .SETN(_0119_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1165_ (.D(_0261_),
    .SETN(_0120_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1166_ (.D(_0262_),
    .SETN(_0121_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1167_ (.D(_0263_),
    .SETN(_0122_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1168_ (.D(_0264_),
    .SETN(_0123_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1169_ (.D(_0265_),
    .SETN(_0124_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1170_ (.D(_0266_),
    .SETN(_0125_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1171_ (.D(_0267_),
    .SETN(_0126_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1172_ (.D(_0268_),
    .SETN(_0127_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1173_ (.D(_0269_),
    .SETN(_0128_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1174_ (.D(_0270_),
    .SETN(_0129_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1175_ (.D(_0271_),
    .SETN(_0130_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1176_ (.D(_0272_),
    .SETN(_0131_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1177_ (.D(_0273_),
    .SETN(_0132_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1178_ (.D(_0274_),
    .SETN(_0133_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1179_ (.D(_0275_),
    .SETN(_0134_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1180_ (.D(_0276_),
    .SETN(_0135_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1181_ (.D(_0277_),
    .SETN(_0136_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1182_ (.D(_0278_),
    .SETN(_0137_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1183_ (.D(_0279_),
    .SETN(_0138_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1184_ (.D(_0280_),
    .SETN(_0139_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1185_ (.D(_0281_),
    .SETN(_0140_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1186_ (.D(_0282_),
    .SETN(_0141_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1187_ (.D(_0283_),
    .SETN(_0142_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1188_ (.D(_0284_),
    .SETN(_0143_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1189_ (.D(_0285_),
    .SETN(_0144_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1190_ (.D(_0286_),
    .SETN(_0145_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1191_ (.D(_0287_),
    .SETN(_0146_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1192_ (.D(_0288_),
    .SETN(_0147_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(preset_n_reg));
 efuse_array_64x32 \efuse_gen_depth[0].efuse_array  (.PRESET_N(preset_n),
    .SENSE(sense),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[31] ,
    \col_prog_n[30] ,
    \col_prog_n[29] ,
    \col_prog_n[28] ,
    \col_prog_n[27] ,
    \col_prog_n[26] ,
    \col_prog_n[25] ,
    \col_prog_n[24] ,
    \col_prog_n[23] ,
    \col_prog_n[22] ,
    \col_prog_n[21] ,
    \col_prog_n[20] ,
    \col_prog_n[19] ,
    \col_prog_n[18] ,
    \col_prog_n[17] ,
    \col_prog_n[16] ,
    \col_prog_n[15] ,
    \col_prog_n[14] ,
    \col_prog_n[13] ,
    \col_prog_n[12] ,
    \col_prog_n[11] ,
    \col_prog_n[10] ,
    \col_prog_n[9] ,
    \col_prog_n[8] ,
    \col_prog_n[7] ,
    \col_prog_n[6] ,
    \col_prog_n[5] ,
    \col_prog_n[4] ,
    \col_prog_n[3] ,
    \col_prog_n[2] ,
    \col_prog_n[1] ,
    \col_prog_n[0] }),
    .OUT({\efuse_out[31] ,
    \efuse_out[30] ,
    \efuse_out[29] ,
    \efuse_out[28] ,
    \efuse_out[27] ,
    \efuse_out[26] ,
    \efuse_out[25] ,
    \efuse_out[24] ,
    \efuse_out[23] ,
    \efuse_out[22] ,
    \efuse_out[21] ,
    \efuse_out[20] ,
    \efuse_out[19] ,
    \efuse_out[18] ,
    \efuse_out[17] ,
    \efuse_out[16] ,
    \efuse_out[15] ,
    \efuse_out[14] ,
    \efuse_out[13] ,
    \efuse_out[12] ,
    \efuse_out[11] ,
    \efuse_out[10] ,
    \efuse_out[9] ,
    \efuse_out[8] ,
    \efuse_out[7] ,
    \efuse_out[6] ,
    \efuse_out[5] ,
    \efuse_out[4] ,
    \efuse_out[3] ,
    \efuse_out[2] ,
    \efuse_out[1] ,
    \efuse_out[0] }));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[0].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[0] ),
    .S(write_enable_i),
    .Z(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[10].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[10] ),
    .S(write_enable_i),
    .Z(\col_prog_n[10] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[11].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[11] ),
    .S(write_enable_i),
    .Z(\col_prog_n[11] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[12].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[12] ),
    .S(write_enable_i),
    .Z(\col_prog_n[12] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[13].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[13] ),
    .S(write_enable_i),
    .Z(\col_prog_n[13] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[14].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[14] ),
    .S(write_enable_i),
    .Z(\col_prog_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[15].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[15] ),
    .S(write_enable_i),
    .Z(\col_prog_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[16].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[16] ),
    .S(write_enable_i),
    .Z(\col_prog_n[16] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[17].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[17] ),
    .S(write_enable_i),
    .Z(\col_prog_n[17] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[18].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[18] ),
    .S(write_enable_i),
    .Z(\col_prog_n[18] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[19].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[19] ),
    .S(write_enable_i),
    .Z(\col_prog_n[19] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[1].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[1] ),
    .S(write_enable_i),
    .Z(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[20].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[20] ),
    .S(write_enable_i),
    .Z(\col_prog_n[20] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[21].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[21] ),
    .S(write_enable_i),
    .Z(\col_prog_n[21] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[22].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[22] ),
    .S(write_enable_i),
    .Z(\col_prog_n[22] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[23].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[23] ),
    .S(write_enable_i),
    .Z(\col_prog_n[23] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[24].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[24] ),
    .S(write_enable_i),
    .Z(\col_prog_n[24] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[25].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[25] ),
    .S(write_enable_i),
    .Z(\col_prog_n[25] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[26].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[26] ),
    .S(write_enable_i),
    .Z(\col_prog_n[26] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[27].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[27] ),
    .S(write_enable_i),
    .Z(\col_prog_n[27] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[28].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[28] ),
    .S(write_enable_i),
    .Z(\col_prog_n[28] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[29].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[29] ),
    .S(write_enable_i),
    .Z(\col_prog_n[29] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[2].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[2] ),
    .S(write_enable_i),
    .Z(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[30].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[30] ),
    .S(write_enable_i),
    .Z(\col_prog_n[30] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[31].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[31] ),
    .S(write_enable_i),
    .Z(\col_prog_n[31] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[3].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[3] ),
    .S(write_enable_i),
    .Z(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[4].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[4] ),
    .S(write_enable_i),
    .Z(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[5].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[5] ),
    .S(write_enable_i),
    .Z(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[6].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[6] ),
    .S(write_enable_i),
    .Z(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[7].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[7] ),
    .S(write_enable_i),
    .Z(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[8].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[8] ),
    .S(write_enable_i),
    .Z(\col_prog_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[9].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[9] ),
    .S(write_enable_i),
    .Z(\col_prog_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[0].bitsel_buf_keep_cell  (.I(\bit_sel_reg[0] ),
    .Z(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[10].bitsel_buf_keep_cell  (.I(\bit_sel_reg[10] ),
    .Z(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[11].bitsel_buf_keep_cell  (.I(\bit_sel_reg[11] ),
    .Z(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[12].bitsel_buf_keep_cell  (.I(\bit_sel_reg[12] ),
    .Z(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[13].bitsel_buf_keep_cell  (.I(\bit_sel_reg[13] ),
    .Z(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[14].bitsel_buf_keep_cell  (.I(\bit_sel_reg[14] ),
    .Z(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[15].bitsel_buf_keep_cell  (.I(\bit_sel_reg[15] ),
    .Z(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[16].bitsel_buf_keep_cell  (.I(\bit_sel_reg[16] ),
    .Z(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[17].bitsel_buf_keep_cell  (.I(\bit_sel_reg[17] ),
    .Z(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[18].bitsel_buf_keep_cell  (.I(\bit_sel_reg[18] ),
    .Z(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[19].bitsel_buf_keep_cell  (.I(\bit_sel_reg[19] ),
    .Z(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[1].bitsel_buf_keep_cell  (.I(\bit_sel_reg[1] ),
    .Z(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[20].bitsel_buf_keep_cell  (.I(\bit_sel_reg[20] ),
    .Z(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[21].bitsel_buf_keep_cell  (.I(\bit_sel_reg[21] ),
    .Z(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[22].bitsel_buf_keep_cell  (.I(\bit_sel_reg[22] ),
    .Z(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[23].bitsel_buf_keep_cell  (.I(\bit_sel_reg[23] ),
    .Z(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[24].bitsel_buf_keep_cell  (.I(\bit_sel_reg[24] ),
    .Z(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[25].bitsel_buf_keep_cell  (.I(\bit_sel_reg[25] ),
    .Z(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[26].bitsel_buf_keep_cell  (.I(\bit_sel_reg[26] ),
    .Z(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[27].bitsel_buf_keep_cell  (.I(\bit_sel_reg[27] ),
    .Z(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[28].bitsel_buf_keep_cell  (.I(\bit_sel_reg[28] ),
    .Z(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[29].bitsel_buf_keep_cell  (.I(\bit_sel_reg[29] ),
    .Z(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[2].bitsel_buf_keep_cell  (.I(\bit_sel_reg[2] ),
    .Z(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[30].bitsel_buf_keep_cell  (.I(\bit_sel_reg[30] ),
    .Z(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[31].bitsel_buf_keep_cell  (.I(\bit_sel_reg[31] ),
    .Z(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[32].bitsel_buf_keep_cell  (.I(\bit_sel_reg[32] ),
    .Z(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[33].bitsel_buf_keep_cell  (.I(\bit_sel_reg[33] ),
    .Z(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[34].bitsel_buf_keep_cell  (.I(\bit_sel_reg[34] ),
    .Z(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[35].bitsel_buf_keep_cell  (.I(\bit_sel_reg[35] ),
    .Z(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[36].bitsel_buf_keep_cell  (.I(\bit_sel_reg[36] ),
    .Z(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[37].bitsel_buf_keep_cell  (.I(\bit_sel_reg[37] ),
    .Z(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[38].bitsel_buf_keep_cell  (.I(\bit_sel_reg[38] ),
    .Z(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[39].bitsel_buf_keep_cell  (.I(\bit_sel_reg[39] ),
    .Z(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[3].bitsel_buf_keep_cell  (.I(\bit_sel_reg[3] ),
    .Z(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[40].bitsel_buf_keep_cell  (.I(\bit_sel_reg[40] ),
    .Z(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[41].bitsel_buf_keep_cell  (.I(\bit_sel_reg[41] ),
    .Z(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[42].bitsel_buf_keep_cell  (.I(\bit_sel_reg[42] ),
    .Z(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[43].bitsel_buf_keep_cell  (.I(\bit_sel_reg[43] ),
    .Z(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[44].bitsel_buf_keep_cell  (.I(\bit_sel_reg[44] ),
    .Z(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[45].bitsel_buf_keep_cell  (.I(\bit_sel_reg[45] ),
    .Z(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[46].bitsel_buf_keep_cell  (.I(\bit_sel_reg[46] ),
    .Z(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[47].bitsel_buf_keep_cell  (.I(\bit_sel_reg[47] ),
    .Z(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[48].bitsel_buf_keep_cell  (.I(\bit_sel_reg[48] ),
    .Z(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[49].bitsel_buf_keep_cell  (.I(\bit_sel_reg[49] ),
    .Z(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[4].bitsel_buf_keep_cell  (.I(\bit_sel_reg[4] ),
    .Z(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[50].bitsel_buf_keep_cell  (.I(\bit_sel_reg[50] ),
    .Z(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[51].bitsel_buf_keep_cell  (.I(\bit_sel_reg[51] ),
    .Z(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[52].bitsel_buf_keep_cell  (.I(\bit_sel_reg[52] ),
    .Z(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[53].bitsel_buf_keep_cell  (.I(\bit_sel_reg[53] ),
    .Z(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[54].bitsel_buf_keep_cell  (.I(\bit_sel_reg[54] ),
    .Z(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[55].bitsel_buf_keep_cell  (.I(\bit_sel_reg[55] ),
    .Z(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[56].bitsel_buf_keep_cell  (.I(\bit_sel_reg[56] ),
    .Z(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[57].bitsel_buf_keep_cell  (.I(\bit_sel_reg[57] ),
    .Z(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[58].bitsel_buf_keep_cell  (.I(\bit_sel_reg[58] ),
    .Z(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[59].bitsel_buf_keep_cell  (.I(\bit_sel_reg[59] ),
    .Z(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[5].bitsel_buf_keep_cell  (.I(\bit_sel_reg[5] ),
    .Z(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[60].bitsel_buf_keep_cell  (.I(\bit_sel_reg[60] ),
    .Z(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[61].bitsel_buf_keep_cell  (.I(\bit_sel_reg[61] ),
    .Z(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[62].bitsel_buf_keep_cell  (.I(\bit_sel_reg[62] ),
    .Z(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[63].bitsel_buf_keep_cell  (.I(\bit_sel_reg[63] ),
    .Z(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[6].bitsel_buf_keep_cell  (.I(\bit_sel_reg[6] ),
    .Z(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[7].bitsel_buf_keep_cell  (.I(\bit_sel_reg[7] ),
    .Z(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[8].bitsel_buf_keep_cell  (.I(\bit_sel_reg[8] ),
    .Z(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[9].bitsel_buf_keep_cell  (.I(\bit_sel_reg[9] ),
    .Z(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].preset_buf_keep_cell  (.I(preset_n_reg),
    .Z(preset_n));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].sense_buf_keep_cell  (.I(sense_del),
    .Z(sense));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[0].sense_dly_keep_cell  (.I(sense_reg),
    .Z(sense_del));
 gf180mcu_fd_sc_mcu7t5v0__tieh tie_keep_cell (.Z(one));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Left_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Left_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Left_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Left_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Left_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Left_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Left_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Left_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Left_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Left_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Left_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Left_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Left_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Left_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Left_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Left_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_2_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_2_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_2_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_2_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_2_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_2_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_2_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_2_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_2_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_2_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_2_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_2_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_2_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_2_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_2_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_2_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_2_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_2_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_2_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_2_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_2_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_2_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_2_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_2_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_2_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_2_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_2_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_2_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_2_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_2_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_2_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_2_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_2_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_2_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_2_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_2_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_2_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_2_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_2_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_2_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_2_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_2_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_2_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_2_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_2_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_2_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_2_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_2_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_2_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_2_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_2_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_2_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_2_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_2_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_2_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_2_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_2_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_2_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_2_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_2_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_2_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_2_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_2_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_2_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_2_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_2_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_2_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_2_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_2_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_2_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_2_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_2_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_2_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_2_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_2_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_2_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_2_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_2_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_2_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_2_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_2_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_2_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_2_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_2_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_2_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_2_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_2_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_2_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_2_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_2_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_2_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_2_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_2_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_2_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_2_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_2_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_2_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_2_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_2_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_2_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_2_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_2_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_2_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_2_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_2_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_2_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_2_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_2_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_2_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_2_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_2_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_2_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_2_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_2_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_2_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_2_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_2_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_2_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_2_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_2_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_2_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_2_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_2_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_2_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_2_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_2_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_2_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_2_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_2_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_2_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_2_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_2_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_2_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_2_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_2_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_2_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_2_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_2_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_2_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_2_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_2_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_2_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_2_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Right_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Right_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Right_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Right_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Right_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Right_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Right_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Right_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Right_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Right_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Right_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Right_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Right_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Right_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Right_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Right_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Right_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Right_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Right_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Right_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Right_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Right_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Right_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Right_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Right_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Right_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Right_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Right_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Right_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Right_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Right_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Right_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Right_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Right_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Right_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Right_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Right_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Right_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Right_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Right_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Right_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Right_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Right_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Right_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Right_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Right_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Right_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Right_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Right_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Right_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Right_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Right_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Right_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Right_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Right_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Right_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Right_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Right_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Right_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Right_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Right_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Right_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Right_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Right_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Right_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Right_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Right_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Right_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Right_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Right_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Right_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Right_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Right_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Right_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Right_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Right_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Right_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Right_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Right_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Right_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Right_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Right_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Right_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Right_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Right_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Right_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Right_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Right_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Right_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Right_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Right_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Right_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Right_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Right_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Right_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Right_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Right_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Right_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Right_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Right_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Right_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Right_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Right_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Right_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Right_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Right_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Right_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Right_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Right_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Right_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Right_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Right_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Right_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Right_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Right_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_2_Right_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_2_Right_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_2_Right_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_2_Right_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_2_Right_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_2_Right_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_2_Right_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_2_Right_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_2_Right_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_2_Right_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_2_Right_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_2_Right_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_2_Right_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_2_Right_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_2_Right_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_2_Right_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_2_Right_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_2_Right_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_2_Right_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_2_Right_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_2_Right_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_2_Right_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_2_Right_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_2_Right_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_2_Right_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_2_Right_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_2_Right_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_2_Right_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_2_Right_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_2_Right_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_2_Right_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_2_Right_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_2_Right_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_2_Right_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_2_Right_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_2_Right_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_2_Right_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_2_Right_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_2_Right_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_2_Right_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_2_Right_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_2_Right_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_2_Right_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_2_Right_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_2_Right_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_2_Right_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_2_Right_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_2_Right_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_2_Right_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_2_Right_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_2_Right_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_2_Right_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_2_Right_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_2_Right_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_2_Right_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_2_Right_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_2_Right_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_2_Right_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_2_Right_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_2_Right_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_2_Right_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_2_Right_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_2_Right_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_2_Right_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_2_Right_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_2_Right_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_2_Right_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_2_Right_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_2_Right_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_2_Right_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_2_Right_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_2_Right_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_2_Right_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_2_Right_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_2_Right_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_2_Right_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_2_Right_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_2_Right_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_2_Right_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_2_Right_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_2_Right_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_2_Right_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_2_Right_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_2_Right_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_2_Right_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_2_Right_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_2_Right_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_2_Right_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_2_Right_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_2_Right_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_2_Right_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_2_Right_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_2_Right_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_2_Right_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_2_Right_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_2_Right_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_2_Right_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_2_Right_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_2_Right_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_2_Right_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_2_Right_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_2_Right_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_2_Right_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_2_Right_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_2_Right_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_2_Right_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_2_Right_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_2_Right_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_2_Right_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_2_Right_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_2_Right_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_2_Right_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_2_Right_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_2_Right_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_2_Right_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_2_Right_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_2_Right_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_2_Right_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_2_Right_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_2_Right_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_2_Right_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_2_Right_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_2_Right_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_2_Right_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_2_Right_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_2_Right_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_2_Right_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_2_Right_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_2_Right_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_2_Right_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_2_Right_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_2_Right_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_2_Right_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_2_Right_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_2_Right_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_2_Right_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_2_Right_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_2_Right_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_2_Right_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_2_Right_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_2_Right_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_2_Right_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_2_Right_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Right_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Right_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Right_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Right_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Right_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Left_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Left_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Left_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Left_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_2_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_2_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_2_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_2_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_2_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_2_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_2_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_2_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_2_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_2_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_2_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_2_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_2_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_2_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_2_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_2_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_2_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_2_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_2_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_2_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_2_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_2_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_2_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_2_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_2_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_2_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_2_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_2_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_2_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_2_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_2_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_2_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_2_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_2_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_2_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_2_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_2_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_2_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_2_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_844 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(wb_adr_i[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(wb_adr_i[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(wb_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(wb_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(wb_adr_i[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(wb_adr_i[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(wb_cyc_i),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(wb_dat_i[0]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(wb_dat_i[10]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(wb_dat_i[11]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(wb_dat_i[12]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(wb_dat_i[13]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(wb_dat_i[14]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(wb_dat_i[15]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(wb_dat_i[16]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(wb_dat_i[17]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(wb_dat_i[18]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(wb_dat_i[19]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(wb_dat_i[1]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(wb_dat_i[20]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(wb_dat_i[21]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(wb_dat_i[22]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(wb_dat_i[23]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(wb_dat_i[24]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(wb_dat_i[25]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(wb_dat_i[26]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(wb_dat_i[27]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(wb_dat_i[28]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(wb_dat_i[29]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(wb_dat_i[2]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(wb_dat_i[30]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(wb_dat_i[31]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(wb_dat_i[3]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(wb_dat_i[4]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(wb_dat_i[5]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(wb_dat_i[6]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(wb_dat_i[7]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(wb_dat_i[8]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(wb_dat_i[9]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(wb_rst_i),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(wb_sel_i[0]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(wb_sel_i[1]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(wb_sel_i[2]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(wb_sel_i[3]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input45 (.I(wb_stb_i),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input46 (.I(wb_we_i),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output47 (.I(net47),
    .Z(wb_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output48 (.I(net48),
    .Z(wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output49 (.I(net49),
    .Z(wb_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output50 (.I(net50),
    .Z(wb_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output51 (.I(net51),
    .Z(wb_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output52 (.I(net52),
    .Z(wb_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output53 (.I(net53),
    .Z(wb_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output54 (.I(net54),
    .Z(wb_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output55 (.I(net55),
    .Z(wb_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output56 (.I(net56),
    .Z(wb_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output57 (.I(net57),
    .Z(wb_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output58 (.I(net58),
    .Z(wb_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output59 (.I(net59),
    .Z(wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output60 (.I(net60),
    .Z(wb_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output61 (.I(net61),
    .Z(wb_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output62 (.I(net62),
    .Z(wb_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output63 (.I(net63),
    .Z(wb_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output64 (.I(net64),
    .Z(wb_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output65 (.I(net65),
    .Z(wb_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output66 (.I(net66),
    .Z(wb_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output67 (.I(net67),
    .Z(wb_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output68 (.I(net68),
    .Z(wb_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output69 (.I(net69),
    .Z(wb_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output70 (.I(net70),
    .Z(wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output71 (.I(net71),
    .Z(wb_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output72 (.I(net72),
    .Z(wb_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output73 (.I(net73),
    .Z(wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output74 (.I(net74),
    .Z(wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output75 (.I(net75),
    .Z(wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output76 (.I(net76),
    .Z(wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output77 (.I(net77),
    .Z(wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output78 (.I(net78),
    .Z(wb_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output79 (.I(net79),
    .Z(wb_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap81 (.I(_0467_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap83 (.I(_0391_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire84 (.I(_0351_),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap85 (.I(_0499_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap87 (.I(_0384_),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew88 (.I(_0291_),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap90 (.I(\state[1] ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew92 (.I(net40),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload0 (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload1 (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload2 (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload3 (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload4 (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload5 (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload6 (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload7 (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_326 ();
endmodule
