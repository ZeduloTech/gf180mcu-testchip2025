module efuse_wb_mem_32x8 (wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rst_i,
    wb_sel_i,
    wb_stb_i,
    wb_we_i,
    write_enable_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o);
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rst_i;
 input wb_sel_i;
 input wb_stb_i;
 input wb_we_i;
 input write_enable_i;
 input [4:0] wb_adr_i;
 input [7:0] wb_dat_i;
 output [7:0] wb_dat_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire \bit_sel[0] ;
 wire \bit_sel[10] ;
 wire \bit_sel[11] ;
 wire \bit_sel[12] ;
 wire \bit_sel[13] ;
 wire \bit_sel[14] ;
 wire \bit_sel[15] ;
 wire \bit_sel[16] ;
 wire \bit_sel[17] ;
 wire \bit_sel[18] ;
 wire \bit_sel[19] ;
 wire \bit_sel[1] ;
 wire \bit_sel[20] ;
 wire \bit_sel[21] ;
 wire \bit_sel[22] ;
 wire \bit_sel[23] ;
 wire \bit_sel[24] ;
 wire \bit_sel[25] ;
 wire \bit_sel[26] ;
 wire \bit_sel[27] ;
 wire \bit_sel[28] ;
 wire \bit_sel[29] ;
 wire \bit_sel[2] ;
 wire \bit_sel[30] ;
 wire \bit_sel[31] ;
 wire \bit_sel[3] ;
 wire \bit_sel[4] ;
 wire \bit_sel[5] ;
 wire \bit_sel[6] ;
 wire \bit_sel[7] ;
 wire \bit_sel[8] ;
 wire \bit_sel[9] ;
 wire \bit_sel_reg[0] ;
 wire \bit_sel_reg[10] ;
 wire \bit_sel_reg[11] ;
 wire \bit_sel_reg[12] ;
 wire \bit_sel_reg[13] ;
 wire \bit_sel_reg[14] ;
 wire \bit_sel_reg[15] ;
 wire \bit_sel_reg[16] ;
 wire \bit_sel_reg[17] ;
 wire \bit_sel_reg[18] ;
 wire \bit_sel_reg[19] ;
 wire \bit_sel_reg[1] ;
 wire \bit_sel_reg[20] ;
 wire \bit_sel_reg[21] ;
 wire \bit_sel_reg[22] ;
 wire \bit_sel_reg[23] ;
 wire \bit_sel_reg[24] ;
 wire \bit_sel_reg[25] ;
 wire \bit_sel_reg[26] ;
 wire \bit_sel_reg[27] ;
 wire \bit_sel_reg[28] ;
 wire \bit_sel_reg[29] ;
 wire \bit_sel_reg[2] ;
 wire \bit_sel_reg[30] ;
 wire \bit_sel_reg[31] ;
 wire \bit_sel_reg[3] ;
 wire \bit_sel_reg[4] ;
 wire \bit_sel_reg[5] ;
 wire \bit_sel_reg[6] ;
 wire \bit_sel_reg[7] ;
 wire \bit_sel_reg[8] ;
 wire \bit_sel_reg[9] ;
 wire \col_prog_n[0] ;
 wire \col_prog_n[1] ;
 wire \col_prog_n[2] ;
 wire \col_prog_n[3] ;
 wire \col_prog_n[4] ;
 wire \col_prog_n[5] ;
 wire \col_prog_n[6] ;
 wire \col_prog_n[7] ;
 wire \col_prog_n_reg[0] ;
 wire \col_prog_n_reg[1] ;
 wire \col_prog_n_reg[2] ;
 wire \col_prog_n_reg[3] ;
 wire \col_prog_n_reg[4] ;
 wire \col_prog_n_reg[5] ;
 wire \col_prog_n_reg[6] ;
 wire \col_prog_n_reg[7] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \efuse_out[0] ;
 wire \efuse_out[1] ;
 wire \efuse_out[2] ;
 wire \efuse_out[3] ;
 wire \efuse_out[4] ;
 wire \efuse_out[5] ;
 wire \efuse_out[6] ;
 wire \efuse_out[7] ;
 wire one;
 wire preset_n;
 wire preset_n_reg;
 wire sense;
 wire sense_del;
 wire sense_reg;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _259_ (.I(preset_n_reg),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _260_ (.I(\col_prog_n_reg[7] ),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _261_ (.I(\state[3] ),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _262_ (.I(\col_prog_n_reg[6] ),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _263_ (.I(\col_prog_n_reg[5] ),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _264_ (.I(\col_prog_n_reg[4] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _265_ (.I(\col_prog_n_reg[3] ),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _266_ (.I(\col_prog_n_reg[2] ),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _267_ (.I(\col_prog_n_reg[1] ),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _268_ (.I(\col_prog_n_reg[0] ),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _269_ (.I(\counter[9] ),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _270_ (.I(\counter[8] ),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _271_ (.I(\counter[7] ),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _272_ (.I(\counter[6] ),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _273_ (.I(\counter[5] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _274_ (.I(\counter[4] ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _275_ (.I(\counter[3] ),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _276_ (.I(\counter[2] ),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _277_ (.I(\counter[1] ),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _278_ (.I(\state[1] ),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _279_ (.I(\state[0] ),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _280_ (.I(net5),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _281_ (.I(net1),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _282_ (.I(net2),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _283_ (.I(net3),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _284_ (.I(net4),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _285_ (.I(net15),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _286_ (.A1(net6),
    .A2(net17),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _287_ (.A1(\state[0] ),
    .A2(net18),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _288_ (.A1(net19),
    .A2(_155_),
    .B(\state[0] ),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _289_ (.A1(net19),
    .A2(net18),
    .A3(_155_),
    .B(\state[0] ),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _290_ (.A1(\state[2] ),
    .A2(_158_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _291_ (.A1(net19),
    .A2(_149_),
    .A3(net18),
    .A4(_155_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _292_ (.A1(_129_),
    .A2(_000_),
    .B(_159_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _293_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .A4(\counter[0] ),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _294_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .A3(\counter[5] ),
    .A4(\counter[4] ),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _295_ (.A1(_140_),
    .A2(_160_),
    .A3(_161_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _296_ (.A1(_140_),
    .A2(_160_),
    .A3(_161_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _297_ (.A1(_131_),
    .A2(_162_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _298_ (.A1(_139_),
    .A2(_140_),
    .A3(_160_),
    .A4(_161_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _299_ (.A1(\state[3] ),
    .A2(_165_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _300_ (.A1(net16),
    .A2(net14),
    .Z(_167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _301_ (.A1(_130_),
    .A2(_131_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _302_ (.A1(net16),
    .A2(net13),
    .Z(_168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _303_ (.A1(_131_),
    .A2(_132_),
    .B1(_166_),
    .B2(_168_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _304_ (.A1(net16),
    .A2(net12),
    .Z(_169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _305_ (.A1(_131_),
    .A2(_133_),
    .B1(_166_),
    .B2(_169_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _306_ (.A1(net16),
    .A2(net11),
    .Z(_170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _307_ (.A1(_131_),
    .A2(_134_),
    .B1(_166_),
    .B2(_170_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _308_ (.A1(net16),
    .A2(net10),
    .Z(_171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _309_ (.A1(_131_),
    .A2(_135_),
    .B1(_166_),
    .B2(_171_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _310_ (.A1(net16),
    .A2(net9),
    .Z(_172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _311_ (.A1(_131_),
    .A2(_136_),
    .B1(_166_),
    .B2(_172_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _312_ (.A1(net16),
    .A2(net8),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _313_ (.A1(_131_),
    .A2(_137_),
    .B1(_166_),
    .B2(_173_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _314_ (.A1(net16),
    .A2(net7),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _315_ (.A1(_131_),
    .A2(_138_),
    .B1(_166_),
    .B2(_174_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _316_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _317_ (.A1(\bit_sel_reg[31] ),
    .A2(_175_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _318_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _319_ (.A1(_154_),
    .A2(_177_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _320_ (.A1(net19),
    .A2(_155_),
    .A3(_156_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _321_ (.A1(net19),
    .A2(_155_),
    .A3(_156_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _322_ (.A1(\state[2] ),
    .A2(_179_),
    .B(net5),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _323_ (.A1(_178_),
    .A2(net29),
    .B(_176_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _324_ (.A1(\bit_sel_reg[30] ),
    .A2(_175_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _325_ (.A1(_151_),
    .A2(net2),
    .A3(net3),
    .A4(net4),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _326_ (.A1(net29),
    .A2(_183_),
    .B(_182_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _327_ (.A1(\bit_sel_reg[29] ),
    .A2(_175_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _328_ (.A1(net1),
    .A2(_152_),
    .A3(net3),
    .A4(net4),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _329_ (.A1(net29),
    .A2(_185_),
    .B(_184_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _330_ (.A1(\bit_sel_reg[28] ),
    .A2(net30),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _331_ (.A1(net1),
    .A2(net2),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _332_ (.A1(net3),
    .A2(net4),
    .A3(_187_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _333_ (.A1(net29),
    .A2(_188_),
    .B(_186_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _334_ (.A1(\bit_sel_reg[27] ),
    .A2(_175_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _335_ (.A1(net1),
    .A2(net2),
    .A3(_153_),
    .A4(net4),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _336_ (.A1(_181_),
    .A2(_190_),
    .B(_189_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _337_ (.A1(\bit_sel_reg[26] ),
    .A2(net30),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _338_ (.A1(net1),
    .A2(_152_),
    .A3(net3),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _339_ (.A1(net4),
    .A2(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _340_ (.A1(net29),
    .A2(_193_),
    .B(_191_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _341_ (.A1(\bit_sel_reg[25] ),
    .A2(net30),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _342_ (.A1(_151_),
    .A2(net2),
    .A3(net3),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _343_ (.A1(net4),
    .A2(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _344_ (.A1(net29),
    .A2(_196_),
    .B(_194_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _345_ (.A1(\bit_sel_reg[24] ),
    .A2(net30),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _346_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _347_ (.A1(net4),
    .A2(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _348_ (.A1(net29),
    .A2(_199_),
    .B(_197_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _349_ (.A1(\bit_sel_reg[23] ),
    .A2(_175_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _350_ (.A1(net4),
    .A2(_177_),
    .A3(net29),
    .B(_200_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _351_ (.A1(\bit_sel_reg[22] ),
    .A2(_175_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _352_ (.A1(_151_),
    .A2(net2),
    .A3(net3),
    .A4(_154_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _353_ (.A1(net29),
    .A2(_202_),
    .B(_201_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _354_ (.A1(\bit_sel_reg[21] ),
    .A2(net30),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _355_ (.A1(net1),
    .A2(_152_),
    .A3(net3),
    .A4(_154_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _356_ (.A1(net29),
    .A2(_204_),
    .B(_203_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _357_ (.A1(\bit_sel_reg[20] ),
    .A2(net30),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _358_ (.A1(net3),
    .A2(_154_),
    .A3(_187_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _359_ (.A1(net29),
    .A2(_206_),
    .B(_205_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _360_ (.A1(\bit_sel_reg[19] ),
    .A2(_175_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _361_ (.A1(net1),
    .A2(net2),
    .A3(_153_),
    .A4(_154_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _362_ (.A1(net29),
    .A2(_208_),
    .B(_207_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _363_ (.A1(\bit_sel_reg[18] ),
    .A2(net30),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _364_ (.A1(_154_),
    .A2(_192_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _365_ (.A1(net29),
    .A2(_210_),
    .B(_209_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _366_ (.A1(\bit_sel_reg[17] ),
    .A2(net30),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _367_ (.A1(_154_),
    .A2(_195_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _368_ (.A1(net29),
    .A2(_212_),
    .B(_211_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _369_ (.A1(\bit_sel_reg[16] ),
    .A2(net30),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _370_ (.A1(_154_),
    .A2(_198_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _371_ (.A1(net29),
    .A2(_214_),
    .B(_213_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _372_ (.A1(\bit_sel_reg[15] ),
    .A2(_175_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _373_ (.A1(\state[2] ),
    .A2(_179_),
    .B(_150_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _374_ (.A1(_178_),
    .A2(net28),
    .B(_215_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _375_ (.A1(\bit_sel_reg[14] ),
    .A2(_175_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _376_ (.A1(_183_),
    .A2(net28),
    .B(_217_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _377_ (.A1(\bit_sel_reg[13] ),
    .A2(_175_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _378_ (.A1(_185_),
    .A2(net28),
    .B(_218_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _379_ (.A1(\bit_sel_reg[12] ),
    .A2(net30),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _380_ (.A1(_188_),
    .A2(net28),
    .B(_219_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _381_ (.A1(\bit_sel_reg[11] ),
    .A2(_175_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _382_ (.A1(_190_),
    .A2(_216_),
    .B(_220_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _383_ (.A1(\bit_sel_reg[10] ),
    .A2(net30),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _384_ (.A1(_193_),
    .A2(net28),
    .B(_221_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _385_ (.A1(\bit_sel_reg[9] ),
    .A2(net30),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _386_ (.A1(_196_),
    .A2(net28),
    .B(_222_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _387_ (.A1(\bit_sel_reg[8] ),
    .A2(net30),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _388_ (.A1(_199_),
    .A2(net28),
    .B(_223_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _389_ (.A1(\bit_sel_reg[7] ),
    .A2(_175_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _390_ (.A1(net4),
    .A2(_177_),
    .A3(net28),
    .B(_224_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _391_ (.A1(\bit_sel_reg[6] ),
    .A2(_175_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _392_ (.A1(_202_),
    .A2(net28),
    .B(_225_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _393_ (.A1(\bit_sel_reg[5] ),
    .A2(net30),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _394_ (.A1(_204_),
    .A2(net28),
    .B(_226_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _395_ (.A1(\bit_sel_reg[4] ),
    .A2(net30),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _396_ (.A1(_206_),
    .A2(net28),
    .B(_227_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _397_ (.A1(\bit_sel_reg[3] ),
    .A2(_175_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _398_ (.A1(_208_),
    .A2(_216_),
    .B(_228_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _399_ (.A1(\bit_sel_reg[2] ),
    .A2(net30),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _400_ (.A1(_210_),
    .A2(net28),
    .B(_229_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _401_ (.A1(\bit_sel_reg[1] ),
    .A2(net30),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _402_ (.A1(_212_),
    .A2(net28),
    .B(_230_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _403_ (.A1(\bit_sel_reg[0] ),
    .A2(net30),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _404_ (.A1(_214_),
    .A2(net28),
    .B(_231_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _405_ (.A1(\state[3] ),
    .A2(_149_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _406_ (.A1(net19),
    .A2(_155_),
    .A3(_156_),
    .B1(\state[0] ),
    .B2(_131_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _407_ (.A1(_162_),
    .A2(_233_),
    .Z(_234_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _408_ (.A1(\state[3] ),
    .A2(_180_),
    .B1(_234_),
    .B2(_139_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _409_ (.A1(_160_),
    .A2(_161_),
    .A3(_233_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _410_ (.A1(_131_),
    .A2(\counter[9] ),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _411_ (.A1(\state[3] ),
    .A2(_139_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _412_ (.A1(_162_),
    .A2(_236_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _413_ (.A1(_180_),
    .A2(_232_),
    .B1(_236_),
    .B2(_162_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _414_ (.A1(_163_),
    .A2(_237_),
    .B(_233_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _415_ (.A1(_140_),
    .A2(_235_),
    .B1(_240_),
    .B2(_164_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _416_ (.A1(_144_),
    .A2(_160_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _417_ (.A1(_143_),
    .A2(_144_),
    .A3(_160_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _418_ (.A1(_142_),
    .A2(_143_),
    .A3(_144_),
    .A4(_160_),
    .Z(_243_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _419_ (.A1(_163_),
    .A2(_237_),
    .B1(_243_),
    .B2(_131_),
    .C(_233_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _420_ (.A1(\state[3] ),
    .A2(_165_),
    .A3(_233_),
    .Z(_245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _421_ (.A1(\state[3] ),
    .A2(_165_),
    .A3(_233_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _422_ (.A1(\counter[7] ),
    .A2(_243_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _423_ (.A1(_141_),
    .A2(_244_),
    .B1(_245_),
    .B2(_247_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _424_ (.A1(_180_),
    .A2(_232_),
    .B1(_236_),
    .B2(_162_),
    .C(_242_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _425_ (.A1(_142_),
    .A2(_248_),
    .B(_244_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _426_ (.A1(_180_),
    .A2(_232_),
    .B1(_236_),
    .B2(_162_),
    .C(_241_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _427_ (.A1(\state[3] ),
    .A2(_180_),
    .B1(_240_),
    .B2(_242_),
    .C1(_249_),
    .C2(_143_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _428_ (.A1(_131_),
    .A2(_160_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _429_ (.A1(_180_),
    .A2(_232_),
    .B1(_236_),
    .B2(_162_),
    .C(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _430_ (.A1(_241_),
    .A2(_246_),
    .B1(_251_),
    .B2(_144_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _431_ (.A1(\counter[2] ),
    .A2(\counter[1] ),
    .A3(\counter[0] ),
    .Z(_252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _432_ (.A1(_180_),
    .A2(_232_),
    .B1(_236_),
    .B2(_162_),
    .C(_252_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _433_ (.A1(_240_),
    .A2(_250_),
    .B1(_253_),
    .B2(_145_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _434_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .B(\counter[2] ),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _435_ (.A1(_252_),
    .A2(_254_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _436_ (.A1(_146_),
    .A2(_239_),
    .B1(_246_),
    .B2(_255_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _437_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Z(_256_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _438_ (.A1(_147_),
    .A2(_239_),
    .B1(_246_),
    .B2(_256_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _439_ (.I0(_245_),
    .I1(_240_),
    .S(\counter[0] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _440_ (.A1(\state[3] ),
    .A2(_149_),
    .B(net19),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _441_ (.A1(\state[3] ),
    .A2(_148_),
    .B(_238_),
    .C(_257_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _442_ (.I0(net27),
    .I1(\efuse_out[7] ),
    .S(\state[1] ),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _443_ (.I0(net26),
    .I1(\efuse_out[6] ),
    .S(\state[1] ),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _444_ (.I0(net25),
    .I1(\efuse_out[5] ),
    .S(\state[1] ),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _445_ (.I0(net24),
    .I1(\efuse_out[4] ),
    .S(\state[1] ),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _446_ (.I0(net23),
    .I1(\efuse_out[3] ),
    .S(\state[1] ),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _447_ (.I0(net22),
    .I1(\efuse_out[2] ),
    .S(\state[1] ),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _448_ (.I0(net21),
    .I1(\efuse_out[1] ),
    .S(\state[1] ),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _449_ (.I0(net20),
    .I1(\efuse_out[0] ),
    .S(\state[1] ),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _450_ (.A1(sense_reg),
    .A2(_000_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _451_ (.A1(\state[1] ),
    .A2(_158_),
    .B(_258_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _452_ (.A1(_148_),
    .A2(_157_),
    .A3(_238_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _453_ (.A1(_166_),
    .A2(_179_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _454_ (.I(net15),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _455_ (.I(net15),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _456_ (.I(net15),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _457_ (.I(net15),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _458_ (.I(net15),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _459_ (.I(net15),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _460_ (.I(net15),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _461_ (.I(net15),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _462_ (.I(net15),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _463_ (.I(net15),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _464_ (.I(net15),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _465_ (.I(net15),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _466_ (.I(net15),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _467_ (.I(net15),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _468_ (.I(net15),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _469_ (.I(net15),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _470_ (.I(net15),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _471_ (.I(net15),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _472_ (.I(net15),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _473_ (.I(net15),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _474_ (.I(net15),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _475_ (.I(net15),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _476_ (.I(net15),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _477_ (.I(net15),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _478_ (.I(net15),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _479_ (.I(net15),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _480_ (.I(net15),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _481_ (.I(net15),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _482_ (.I(net15),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _483_ (.I(net15),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _484_ (.I(net15),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _485_ (.I(net15),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _486_ (.I(net15),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _487_ (.I(net15),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _488_ (.I(net15),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _489_ (.I(net15),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _490_ (.I(net15),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _491_ (.I(net15),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _492_ (.I(net15),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _493_ (.I(net15),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _494_ (.I(net15),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _495_ (.I(net15),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _496_ (.I(net15),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _497_ (.I(net15),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _498_ (.I(net15),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _499_ (.I(net15),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _500_ (.I(net15),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _501_ (.I(net15),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _502_ (.I(net15),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _503_ (.I(net15),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _504_ (.I(net15),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _505_ (.I(net15),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _506_ (.I(net15),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _507_ (.I(net15),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _508_ (.I(net15),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _509_ (.I(net15),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _510_ (.I(net15),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _511_ (.I(net15),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _512_ (.I(net15),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _513_ (.I(net15),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _514_ (.I(net15),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _515_ (.I(net15),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _516_ (.I(net15),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _517_ (.I(net15),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _518_ (.D(_068_),
    .RN(_003_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(sense_reg));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _519_ (.D(_069_),
    .RN(_004_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _520_ (.D(_070_),
    .RN(_005_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _521_ (.D(_071_),
    .RN(_006_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _522_ (.D(_072_),
    .RN(_007_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _523_ (.D(_073_),
    .RN(_008_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _524_ (.D(_074_),
    .RN(_009_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _525_ (.D(_075_),
    .RN(_010_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _526_ (.D(_076_),
    .RN(_011_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _527_ (.D(_077_),
    .RN(_012_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _528_ (.D(_078_),
    .RN(_013_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _529_ (.D(_079_),
    .RN(_014_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _530_ (.D(_080_),
    .RN(_015_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _531_ (.D(_081_),
    .RN(_016_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _532_ (.D(_082_),
    .RN(_017_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _533_ (.D(_083_),
    .RN(_018_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _534_ (.D(_084_),
    .RN(_019_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _535_ (.D(_085_),
    .RN(_020_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _536_ (.D(_086_),
    .RN(_021_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _537_ (.D(_087_),
    .RN(_022_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _538_ (.D(_088_),
    .RN(_023_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _539_ (.D(_089_),
    .RN(_024_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _540_ (.D(_090_),
    .RN(_025_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _541_ (.D(_091_),
    .RN(_026_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _542_ (.D(_092_),
    .RN(_027_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _543_ (.D(_093_),
    .RN(_028_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _544_ (.D(_094_),
    .RN(_029_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _545_ (.D(_095_),
    .RN(_030_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _546_ (.D(_096_),
    .RN(_031_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _547_ (.D(_097_),
    .RN(_032_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _548_ (.D(_098_),
    .RN(_033_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _549_ (.D(_099_),
    .RN(_034_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _550_ (.D(_100_),
    .RN(_035_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _551_ (.D(_101_),
    .RN(_036_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _552_ (.D(_102_),
    .RN(_037_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _553_ (.D(_103_),
    .RN(_038_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _554_ (.D(_104_),
    .RN(_039_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _555_ (.D(_105_),
    .RN(_040_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _556_ (.D(_106_),
    .RN(_041_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _557_ (.D(_107_),
    .RN(_042_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _558_ (.D(_108_),
    .RN(_043_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _559_ (.D(_109_),
    .RN(_044_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _560_ (.D(_110_),
    .RN(_045_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _561_ (.D(_111_),
    .RN(_046_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _562_ (.D(_112_),
    .RN(_047_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _563_ (.D(_113_),
    .RN(_048_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _564_ (.D(_114_),
    .RN(_049_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _565_ (.D(_115_),
    .RN(_050_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\bit_sel_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _566_ (.D(_116_),
    .RN(_051_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _567_ (.D(_117_),
    .RN(_052_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _568_ (.D(_118_),
    .RN(_053_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _569_ (.D(_119_),
    .RN(_054_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _570_ (.D(_120_),
    .SETN(_055_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _571_ (.D(_121_),
    .SETN(_056_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _572_ (.D(_122_),
    .SETN(_057_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _573_ (.D(_123_),
    .SETN(_058_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _574_ (.D(_124_),
    .SETN(_059_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _575_ (.D(_125_),
    .SETN(_060_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _576_ (.D(_126_),
    .SETN(_061_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _577_ (.D(_127_),
    .SETN(_062_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _578_ (.D(_128_),
    .SETN(_063_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(preset_n_reg));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _579_ (.D(_001_),
    .SETN(_064_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _580_ (.D(\state[2] ),
    .RN(_065_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _581_ (.D(_000_),
    .RN(_066_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _582_ (.D(_002_),
    .RN(_067_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\state[3] ));
 efuse_array_32x8 \efuse_gen_depth[0].efuse_array  (.PRESET_N(preset_n),
    .SENSE(sense),
    .BIT_SEL({\bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[7] ,
    \col_prog_n[6] ,
    \col_prog_n[5] ,
    \col_prog_n[4] ,
    \col_prog_n[3] ,
    \col_prog_n[2] ,
    \col_prog_n[1] ,
    \col_prog_n[0] }),
    .OUT({\efuse_out[7] ,
    \efuse_out[6] ,
    \efuse_out[5] ,
    \efuse_out[4] ,
    \efuse_out[3] ,
    \efuse_out[2] ,
    \efuse_out[1] ,
    \efuse_out[0] }));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[0].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[0] ),
    .S(write_enable_i),
    .Z(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[1].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[1] ),
    .S(write_enable_i),
    .Z(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[2].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[2] ),
    .S(write_enable_i),
    .Z(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[3].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[3] ),
    .S(write_enable_i),
    .Z(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[4].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[4] ),
    .S(write_enable_i),
    .Z(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[5].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[5] ),
    .S(write_enable_i),
    .Z(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[6].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[6] ),
    .S(write_enable_i),
    .Z(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[7].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[7] ),
    .S(write_enable_i),
    .Z(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[0].bitsel_buf_keep_cell  (.I(\bit_sel_reg[0] ),
    .Z(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[10].bitsel_buf_keep_cell  (.I(\bit_sel_reg[10] ),
    .Z(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[11].bitsel_buf_keep_cell  (.I(\bit_sel_reg[11] ),
    .Z(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[12].bitsel_buf_keep_cell  (.I(\bit_sel_reg[12] ),
    .Z(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[13].bitsel_buf_keep_cell  (.I(\bit_sel_reg[13] ),
    .Z(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[14].bitsel_buf_keep_cell  (.I(\bit_sel_reg[14] ),
    .Z(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[15].bitsel_buf_keep_cell  (.I(\bit_sel_reg[15] ),
    .Z(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[16].bitsel_buf_keep_cell  (.I(\bit_sel_reg[16] ),
    .Z(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[17].bitsel_buf_keep_cell  (.I(\bit_sel_reg[17] ),
    .Z(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[18].bitsel_buf_keep_cell  (.I(\bit_sel_reg[18] ),
    .Z(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[19].bitsel_buf_keep_cell  (.I(\bit_sel_reg[19] ),
    .Z(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[1].bitsel_buf_keep_cell  (.I(\bit_sel_reg[1] ),
    .Z(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[20].bitsel_buf_keep_cell  (.I(\bit_sel_reg[20] ),
    .Z(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[21].bitsel_buf_keep_cell  (.I(\bit_sel_reg[21] ),
    .Z(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[22].bitsel_buf_keep_cell  (.I(\bit_sel_reg[22] ),
    .Z(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[23].bitsel_buf_keep_cell  (.I(\bit_sel_reg[23] ),
    .Z(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[24].bitsel_buf_keep_cell  (.I(\bit_sel_reg[24] ),
    .Z(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[25].bitsel_buf_keep_cell  (.I(\bit_sel_reg[25] ),
    .Z(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[26].bitsel_buf_keep_cell  (.I(\bit_sel_reg[26] ),
    .Z(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[27].bitsel_buf_keep_cell  (.I(\bit_sel_reg[27] ),
    .Z(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[28].bitsel_buf_keep_cell  (.I(\bit_sel_reg[28] ),
    .Z(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[29].bitsel_buf_keep_cell  (.I(\bit_sel_reg[29] ),
    .Z(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[2].bitsel_buf_keep_cell  (.I(\bit_sel_reg[2] ),
    .Z(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[30].bitsel_buf_keep_cell  (.I(\bit_sel_reg[30] ),
    .Z(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[31].bitsel_buf_keep_cell  (.I(\bit_sel_reg[31] ),
    .Z(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[3].bitsel_buf_keep_cell  (.I(\bit_sel_reg[3] ),
    .Z(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[4].bitsel_buf_keep_cell  (.I(\bit_sel_reg[4] ),
    .Z(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[5].bitsel_buf_keep_cell  (.I(\bit_sel_reg[5] ),
    .Z(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[6].bitsel_buf_keep_cell  (.I(\bit_sel_reg[6] ),
    .Z(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[7].bitsel_buf_keep_cell  (.I(\bit_sel_reg[7] ),
    .Z(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[8].bitsel_buf_keep_cell  (.I(\bit_sel_reg[8] ),
    .Z(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[9].bitsel_buf_keep_cell  (.I(\bit_sel_reg[9] ),
    .Z(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].preset_buf_keep_cell  (.I(preset_n_reg),
    .Z(preset_n));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].sense_buf_keep_cell  (.I(sense_del),
    .Z(sense));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[0].sense_dly_keep_cell  (.I(sense_reg),
    .Z(sense_del));
 gf180mcu_fd_sc_mcu7t5v0__tieh tie_keep_cell (.Z(one));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Left_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Left_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Left_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Left_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Left_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Left_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Left_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Left_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Left_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Left_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Left_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Left_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Left_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Left_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Left_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Left_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_2_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_2_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_2_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_2_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_2_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_2_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_2_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_2_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_2_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(wb_adr_i[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(wb_adr_i[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(wb_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(wb_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(wb_adr_i[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(wb_cyc_i),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(wb_dat_i[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(wb_dat_i[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(wb_dat_i[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(wb_dat_i[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(wb_dat_i[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(wb_dat_i[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(wb_dat_i[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(wb_dat_i[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(wb_rst_i),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(wb_sel_i),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(wb_stb_i),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(wb_we_i),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output19 (.I(net19),
    .Z(wb_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output20 (.I(net20),
    .Z(wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output21 (.I(net21),
    .Z(wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output22 (.I(net22),
    .Z(wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output23 (.I(net23),
    .Z(wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output24 (.I(net24),
    .Z(wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output25 (.I(net25),
    .Z(wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output26 (.I(net26),
    .Z(wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output27 (.I(net27),
    .Z(wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap28 (.I(_216_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire29 (.I(_181_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap30 (.I(_175_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload0 (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload1 (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload2 (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload3 (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload4 (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload5 (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload6 (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_adr_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(wb_adr_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(wb_adr_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(wb_adr_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(wb_adr_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(wb_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(wb_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(wb_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(wb_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wb_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(wb_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(wb_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(wb_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(wb_sel_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(wb_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(wb_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[7].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[6].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[5].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[4].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[3].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[2].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[1].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[0].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[0].prog_disable_keep_cell_Z  (.I(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[0]  (.I(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[0]  (.I(\efuse_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__I1 (.I(\efuse_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[1]  (.I(\efuse_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__I1 (.I(\efuse_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_Z (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__486__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__479__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__467__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_358 ();
endmodule
