VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_wb_mem_128x8
  CLASS BLOCK ;
  FOREIGN efuse_wb_mem_128x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 464.460 BY 365.825 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.080 2.760 6.080 361.800 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 2.760 460.160 4.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 359.800 460.160 361.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 458.160 2.760 460.160 361.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 0.260 15.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 341.385 15.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.280 0.260 65.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 0.260 115.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 340.760 115.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 0.260 165.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.280 0.260 215.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 264.280 0.260 265.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.280 0.260 315.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.280 341.385 315.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.280 0.260 365.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 414.280 0.260 415.880 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 15.960 462.660 17.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 65.960 462.660 67.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 115.960 462.660 117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 165.960 462.660 167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 215.960 462.660 217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 265.960 462.660 267.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 315.960 462.660 317.560 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 1.580 0.260 3.580 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 0.260 462.660 2.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 362.300 462.660 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 460.660 0.260 462.660 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 0.260 19.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 340.740 19.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.580 0.260 69.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 0.260 119.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 340.740 119.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 0.260 169.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.580 0.260 219.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 267.580 0.260 269.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 317.580 0.260 319.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 367.580 0.260 369.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 367.580 340.740 369.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 417.580 0.260 419.180 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 19.260 462.660 20.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 69.260 462.660 70.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 119.260 462.660 120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 169.260 462.660 170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 219.260 462.660 220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 269.260 462.660 270.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 319.260 462.660 320.860 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 365.265 43.120 365.825 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 365.265 101.360 365.825 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 365.265 115.920 365.825 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 365.265 130.480 365.825 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 365.265 145.040 365.825 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 365.265 159.600 365.825 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 365.265 174.160 365.825 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 365.265 188.720 365.825 ;
    END
  END wb_adr_i[6]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 365.265 72.240 365.825 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 365.265 28.560 365.825 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 365.265 203.280 365.825 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 365.265 217.840 365.825 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 365.265 232.400 365.825 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 365.265 246.960 365.825 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 365.265 261.520 365.825 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 365.265 276.080 365.825 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 365.265 290.640 365.825 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 365.265 305.200 365.825 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 365.265 334.320 365.825 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 365.265 348.880 365.825 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 365.265 363.440 365.825 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 365.265 378.000 365.825 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 365.265 392.560 365.825 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 365.265 407.120 365.825 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 365.265 421.680 365.825 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 365.265 436.240 365.825 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 365.265 57.680 365.825 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 365.265 319.760 365.825 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 365.265 14.000 365.825 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 365.265 86.800 365.825 ;
    END
  END wb_we_i
  PIN write_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 35.264000 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 365.265 450.800 365.825 ;
    END
  END write_enable_i
  OBS
      LAYER Nwell ;
        RECT 9.650 11.330 454.590 353.230 ;
      LAYER Metal1 ;
        RECT 10.080 11.460 454.160 353.100 ;
      LAYER Metal2 ;
        RECT 7.980 364.965 13.140 365.685 ;
        RECT 14.300 364.965 27.700 365.685 ;
        RECT 28.860 364.965 42.260 365.685 ;
        RECT 43.420 364.965 56.820 365.685 ;
        RECT 57.980 364.965 71.380 365.685 ;
        RECT 72.540 364.965 85.940 365.685 ;
        RECT 87.100 364.965 100.500 365.685 ;
        RECT 101.660 364.965 115.060 365.685 ;
        RECT 116.220 364.965 129.620 365.685 ;
        RECT 130.780 364.965 144.180 365.685 ;
        RECT 145.340 364.965 158.740 365.685 ;
        RECT 159.900 364.965 173.300 365.685 ;
        RECT 174.460 364.965 187.860 365.685 ;
        RECT 189.020 364.965 202.420 365.685 ;
        RECT 203.580 364.965 216.980 365.685 ;
        RECT 218.140 364.965 231.540 365.685 ;
        RECT 232.700 364.965 246.100 365.685 ;
        RECT 247.260 364.965 260.660 365.685 ;
        RECT 261.820 364.965 275.220 365.685 ;
        RECT 276.380 364.965 289.780 365.685 ;
        RECT 290.940 364.965 304.340 365.685 ;
        RECT 305.500 364.965 318.900 365.685 ;
        RECT 320.060 364.965 333.460 365.685 ;
        RECT 334.620 364.965 348.020 365.685 ;
        RECT 349.180 364.965 362.580 365.685 ;
        RECT 363.740 364.965 377.140 365.685 ;
        RECT 378.300 364.965 391.700 365.685 ;
        RECT 392.860 364.965 406.260 365.685 ;
        RECT 407.420 364.965 420.820 365.685 ;
        RECT 421.980 364.965 435.380 365.685 ;
        RECT 436.540 364.965 449.940 365.685 ;
        RECT 7.980 5.130 450.660 364.965 ;
      LAYER Metal3 ;
        RECT 7.930 5.180 450.710 365.540 ;
      LAYER Metal4 ;
        RECT 10.240 364.600 383.820 365.590 ;
        RECT 10.240 341.085 13.980 364.600 ;
        RECT 16.180 341.085 17.280 364.600 ;
        RECT 10.240 340.440 17.280 341.085 ;
        RECT 19.480 340.440 63.980 364.600 ;
        RECT 10.240 5.130 63.980 340.440 ;
        RECT 66.180 5.130 67.280 364.600 ;
        RECT 69.480 340.460 113.980 364.600 ;
        RECT 116.180 340.460 117.280 364.600 ;
        RECT 69.480 340.440 117.280 340.460 ;
        RECT 119.480 340.440 163.980 364.600 ;
        RECT 69.480 5.130 163.980 340.440 ;
        RECT 166.180 5.130 167.280 364.600 ;
        RECT 169.480 5.130 213.980 364.600 ;
        RECT 216.180 5.130 217.280 364.600 ;
        RECT 219.480 5.130 263.980 364.600 ;
        RECT 266.180 5.130 267.280 364.600 ;
        RECT 269.480 341.085 313.980 364.600 ;
        RECT 316.180 341.085 317.280 364.600 ;
        RECT 269.480 5.130 317.280 341.085 ;
        RECT 319.480 5.130 363.980 364.600 ;
        RECT 366.180 340.440 367.280 364.600 ;
        RECT 369.480 340.440 383.820 364.600 ;
        RECT 366.180 5.130 383.820 340.440 ;
  END
END efuse_wb_mem_128x8
END LIBRARY

