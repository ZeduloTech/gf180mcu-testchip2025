// Caravel pad assignment

`ifndef _PINOUT_VH
`define _PINOUT_VH

`define NUM_INPUT_PADS  12
`define NUM_BIDIR_PADS  42

`define PAD_CARAVELIO_0 0
`define PAD_GPIO        13
`define PAD_FLASH_CSB   14
`define PAD_FLASH_CLK   15
`define PAD_FLASH_IO0   16
`define PAD_FLASH_IO1   17

`endif
