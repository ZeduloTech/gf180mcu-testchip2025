VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_wb_mem_32x8
  CLASS BLOCK ;
  FOREIGN efuse_wb_mem_32x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 222.730 BY 365.825 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.080 2.760 6.080 361.800 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 2.760 218.240 4.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 359.800 218.240 361.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.240 2.760 218.240 361.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 0.260 15.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 341.385 15.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.280 0.260 65.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 0.260 115.880 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 0.260 165.880 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 15.960 220.740 17.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 65.960 220.740 67.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 115.960 220.740 117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 165.960 220.740 167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 215.960 220.740 217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 265.960 220.740 267.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 315.960 220.740 317.560 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 1.580 0.260 3.580 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 0.260 220.740 2.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 362.300 220.740 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.740 0.260 220.740 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 0.260 19.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 340.740 19.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.580 0.260 69.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 0.260 119.180 364.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 0.260 169.180 364.300 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 19.260 220.740 20.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 69.260 220.740 70.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 119.260 220.740 120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 169.260 220.740 170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 219.260 220.740 220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 269.260 220.740 270.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 319.260 220.740 320.860 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 365.265 30.800 365.825 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 365.265 57.680 365.825 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 365.265 64.400 365.825 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 365.265 71.120 365.825 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 365.265 77.840 365.825 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 365.265 84.560 365.825 ;
    END
  END wb_adr_i[4]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 365.265 44.240 365.825 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 365.265 24.080 365.825 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 365.265 91.280 365.825 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 365.265 98.000 365.825 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 365.265 104.720 365.825 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 365.265 111.440 365.825 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 365.265 118.160 365.825 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 365.265 124.880 365.825 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 365.265 131.600 365.825 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 365.265 138.320 365.825 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 365.265 151.760 365.825 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 365.265 158.480 365.825 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 365.265 165.200 365.825 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 365.265 171.920 365.825 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 365.265 178.640 365.825 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 365.265 185.360 365.825 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 365.265 192.080 365.825 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 365.265 198.800 365.825 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 365.265 37.520 365.825 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 365.265 145.040 365.825 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 365.265 17.360 365.825 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 365.265 50.960 365.825 ;
    END
  END wb_we_i
  PIN write_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 17.632000 ;
    ANTENNADIFFAREA 3.283200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 365.265 205.520 365.825 ;
    END
  END write_enable_i
  OBS
      LAYER Nwell ;
        RECT 9.650 11.330 212.670 353.230 ;
      LAYER Metal1 ;
        RECT 10.080 11.460 212.240 353.100 ;
      LAYER Metal2 ;
        RECT 9.100 364.965 16.500 365.685 ;
        RECT 17.660 364.965 23.220 365.685 ;
        RECT 24.380 364.965 29.940 365.685 ;
        RECT 31.100 364.965 36.660 365.685 ;
        RECT 37.820 364.965 43.380 365.685 ;
        RECT 44.540 364.965 50.100 365.685 ;
        RECT 51.260 364.965 56.820 365.685 ;
        RECT 57.980 364.965 63.540 365.685 ;
        RECT 64.700 364.965 70.260 365.685 ;
        RECT 71.420 364.965 76.980 365.685 ;
        RECT 78.140 364.965 83.700 365.685 ;
        RECT 84.860 364.965 90.420 365.685 ;
        RECT 91.580 364.965 97.140 365.685 ;
        RECT 98.300 364.965 103.860 365.685 ;
        RECT 105.020 364.965 110.580 365.685 ;
        RECT 111.740 364.965 117.300 365.685 ;
        RECT 118.460 364.965 124.020 365.685 ;
        RECT 125.180 364.965 130.740 365.685 ;
        RECT 131.900 364.965 137.460 365.685 ;
        RECT 138.620 364.965 144.180 365.685 ;
        RECT 145.340 364.965 150.900 365.685 ;
        RECT 152.060 364.965 157.620 365.685 ;
        RECT 158.780 364.965 164.340 365.685 ;
        RECT 165.500 364.965 171.060 365.685 ;
        RECT 172.220 364.965 177.780 365.685 ;
        RECT 178.940 364.965 184.500 365.685 ;
        RECT 185.660 364.965 191.220 365.685 ;
        RECT 192.380 364.965 197.940 365.685 ;
        RECT 199.100 364.965 204.660 365.685 ;
        RECT 9.100 11.570 205.380 364.965 ;
      LAYER Metal3 ;
        RECT 10.270 11.620 205.430 364.980 ;
      LAYER Metal4 ;
        RECT 10.240 364.600 161.140 365.030 ;
        RECT 10.240 341.085 13.980 364.600 ;
        RECT 16.180 341.085 17.280 364.600 ;
        RECT 10.240 340.440 17.280 341.085 ;
        RECT 19.480 340.440 63.980 364.600 ;
        RECT 10.240 12.970 63.980 340.440 ;
        RECT 66.180 12.970 67.280 364.600 ;
        RECT 69.480 12.970 113.980 364.600 ;
        RECT 116.180 12.970 117.280 364.600 ;
        RECT 119.480 12.970 161.140 364.600 ;
  END
END efuse_wb_mem_32x8
END LIBRARY

