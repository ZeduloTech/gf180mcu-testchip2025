VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_wb_mem_64x8
  CLASS BLOCK ;
  FOREIGN efuse_wb_mem_64x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 240.000 BY 350.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.080 2.760 6.080 346.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 2.760 235.600 4.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 344.120 235.600 346.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 233.600 2.760 235.600 346.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 0.260 15.880 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.280 0.260 65.880 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 0.260 115.880 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 0.260 165.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 340.760 165.880 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.280 0.260 215.880 348.620 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 15.960 238.100 17.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 65.960 238.100 67.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 115.960 238.100 117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 165.960 238.100 167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 215.960 238.100 217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 265.960 238.100 267.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 315.960 238.100 317.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.600 11.460 226.200 337.420 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 1.580 0.260 3.580 348.620 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 0.260 238.100 2.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 346.620 238.100 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 236.100 0.260 238.100 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 0.260 19.180 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.580 0.260 69.180 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 0.260 119.180 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 0.260 169.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 340.760 169.180 348.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.580 0.260 219.180 348.620 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 19.260 238.100 20.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 69.260 238.100 70.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 119.260 238.100 120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 169.260 238.100 170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 219.260 238.100 220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 269.260 238.100 270.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 319.260 238.100 320.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 226.840 11.460 228.440 337.420 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 349.440 31.920 350.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 349.440 58.800 350.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 349.440 65.520 350.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 349.440 72.240 350.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 349.440 78.960 350.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 349.440 85.680 350.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 349.440 92.400 350.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 349.440 99.120 350.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 349.440 105.840 350.000 ;
    END
  END wb_adr_i[7]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 349.440 45.360 350.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 349.440 25.200 350.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 349.440 112.560 350.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 349.440 119.280 350.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 349.440 126.000 350.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 349.440 132.720 350.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 349.440 139.440 350.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 349.440 146.160 350.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 349.440 152.880 350.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 349.440 159.600 350.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 349.440 166.320 350.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 349.440 173.040 350.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 349.440 179.760 350.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 349.440 186.480 350.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 349.440 193.200 350.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 349.440 199.920 350.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 349.440 206.640 350.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 349.440 213.360 350.000 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 349.440 38.640 350.000 ;
    END
  END wb_rst_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 349.440 18.480 350.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 349.440 52.080 350.000 ;
    END
  END wb_we_i
  PIN write_disable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 17.632000 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 349.440 220.080 350.000 ;
    END
  END write_disable_i
  OBS
      LAYER Nwell ;
        RECT 9.650 11.330 230.030 337.550 ;
      LAYER Metal1 ;
        RECT 10.080 11.460 229.600 337.420 ;
      LAYER Metal2 ;
        RECT 0.140 349.140 17.620 349.860 ;
        RECT 18.780 349.140 24.340 349.860 ;
        RECT 25.500 349.140 31.060 349.860 ;
        RECT 32.220 349.140 37.780 349.860 ;
        RECT 38.940 349.140 44.500 349.860 ;
        RECT 45.660 349.140 51.220 349.860 ;
        RECT 52.380 349.140 57.940 349.860 ;
        RECT 59.100 349.140 64.660 349.860 ;
        RECT 65.820 349.140 71.380 349.860 ;
        RECT 72.540 349.140 78.100 349.860 ;
        RECT 79.260 349.140 84.820 349.860 ;
        RECT 85.980 349.140 91.540 349.860 ;
        RECT 92.700 349.140 98.260 349.860 ;
        RECT 99.420 349.140 104.980 349.860 ;
        RECT 106.140 349.140 111.700 349.860 ;
        RECT 112.860 349.140 118.420 349.860 ;
        RECT 119.580 349.140 125.140 349.860 ;
        RECT 126.300 349.140 131.860 349.860 ;
        RECT 133.020 349.140 138.580 349.860 ;
        RECT 139.740 349.140 145.300 349.860 ;
        RECT 146.460 349.140 152.020 349.860 ;
        RECT 153.180 349.140 158.740 349.860 ;
        RECT 159.900 349.140 165.460 349.860 ;
        RECT 166.620 349.140 172.180 349.860 ;
        RECT 173.340 349.140 178.900 349.860 ;
        RECT 180.060 349.140 185.620 349.860 ;
        RECT 186.780 349.140 192.340 349.860 ;
        RECT 193.500 349.140 199.060 349.860 ;
        RECT 200.220 349.140 205.780 349.860 ;
        RECT 206.940 349.140 212.500 349.860 ;
        RECT 213.660 349.140 219.220 349.860 ;
        RECT 220.380 349.140 232.820 349.860 ;
        RECT 0.140 0.650 232.820 349.140 ;
      LAYER Metal3 ;
        RECT 0.090 0.700 232.870 349.300 ;
      LAYER Metal4 ;
        RECT 0.140 0.650 1.280 343.190 ;
        RECT 6.380 2.460 13.980 343.190 ;
        RECT 3.880 0.650 13.980 2.460 ;
        RECT 16.180 0.650 17.280 343.190 ;
        RECT 19.480 0.650 63.980 343.190 ;
        RECT 66.180 0.650 67.280 343.190 ;
        RECT 69.480 0.650 113.980 343.190 ;
        RECT 116.180 0.650 117.280 343.190 ;
        RECT 119.480 340.460 163.980 343.190 ;
        RECT 166.180 340.460 167.280 343.190 ;
        RECT 169.480 340.460 213.980 343.190 ;
        RECT 119.480 4.740 213.980 340.460 ;
        RECT 119.480 0.650 163.980 4.740 ;
        RECT 166.180 0.650 167.280 4.740 ;
        RECT 169.480 0.650 213.980 4.740 ;
        RECT 216.180 0.650 217.280 343.190 ;
        RECT 219.480 337.720 231.700 343.190 ;
        RECT 219.480 11.160 224.300 337.720 ;
        RECT 226.500 11.160 226.540 337.720 ;
        RECT 228.740 11.160 231.700 337.720 ;
        RECT 219.480 0.650 231.700 11.160 ;
      LAYER Metal5 ;
        RECT 6.780 321.360 231.780 331.870 ;
        RECT 6.780 318.060 231.780 318.760 ;
        RECT 6.780 271.360 231.780 315.460 ;
        RECT 6.780 268.060 231.780 268.760 ;
        RECT 6.780 221.360 231.780 265.460 ;
        RECT 6.780 218.060 231.780 218.760 ;
        RECT 6.780 171.360 231.780 215.460 ;
        RECT 6.780 168.060 231.780 168.760 ;
        RECT 6.780 121.360 231.780 165.460 ;
        RECT 6.780 118.060 231.780 118.760 ;
        RECT 6.780 71.360 231.780 115.460 ;
        RECT 6.780 68.060 231.780 68.760 ;
        RECT 6.780 21.360 231.780 65.460 ;
        RECT 6.780 18.060 231.780 18.760 ;
        RECT 6.780 5.630 231.780 15.460 ;
  END
END efuse_wb_mem_64x8
END LIBRARY

