VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_wb_mem_1024x32
  CLASS BLOCK ;
  FOREIGN efuse_wb_mem_1024x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2856.480 BY 1311.065 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.080 2.760 6.080 1306.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 2.760 2852.480 4.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.080 1304.520 2852.480 1306.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2850.480 2.760 2852.480 1306.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 0.260 15.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.280 1286.625 15.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.280 0.260 65.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 0.260 115.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.280 1285.580 115.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 164.280 0.260 165.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.280 0.260 215.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 264.280 0.260 265.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.280 0.260 315.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.280 1285.580 315.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.280 0.260 365.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 414.280 0.260 415.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 414.280 1285.580 415.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 464.280 0.260 465.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 514.280 0.260 515.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 564.280 0.260 565.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 614.280 0.260 615.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 614.280 1285.580 615.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.280 0.260 665.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 714.280 0.260 715.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 764.280 0.260 765.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 764.280 1285.580 765.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 814.280 0.260 815.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.280 0.260 865.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.280 1286.625 865.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 914.280 0.260 915.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 964.280 0.260 965.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 964.280 1285.580 965.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1014.280 0.260 1015.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1064.280 0.260 1065.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.280 0.260 1115.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.280 1286.625 1115.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1164.280 0.260 1165.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1214.280 0.260 1215.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1214.280 1286.625 1215.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.280 0.260 1265.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1264.280 1286.625 1265.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1314.280 0.260 1315.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1364.280 0.260 1365.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1364.280 1286.625 1365.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1414.280 0.260 1415.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1464.280 0.260 1465.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1514.280 0.260 1515.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1514.280 1285.580 1515.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1564.280 0.260 1565.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1614.280 0.260 1615.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1664.280 0.260 1665.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1714.280 0.260 1715.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1714.280 1285.580 1715.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1764.280 0.260 1765.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1814.280 0.260 1815.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1864.280 0.260 1865.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1864.280 1286.625 1865.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1914.280 0.260 1915.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1964.280 0.260 1965.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2014.280 0.260 2015.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2014.280 1286.625 2015.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2064.280 0.260 2065.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2114.280 0.260 2115.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2114.280 1286.625 2115.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2164.280 0.260 2165.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2164.280 1285.580 2165.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2214.280 0.260 2215.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2264.280 0.260 2265.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2264.280 1285.580 2265.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2314.280 0.260 2315.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2364.280 0.260 2365.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2364.280 1285.580 2365.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2414.280 0.260 2415.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.280 0.260 2465.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.280 1285.580 2465.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2514.280 0.260 2515.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2514.280 1286.625 2515.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2564.280 0.260 2565.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2614.280 0.260 2615.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2614.280 1285.580 2615.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2664.280 0.260 2665.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2714.280 0.260 2715.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2714.280 1285.580 2715.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2764.280 0.260 2765.880 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2814.280 0.260 2815.880 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2814.280 1285.580 2815.880 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 15.960 2854.980 17.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 65.960 2854.980 67.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 115.960 2854.980 117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 165.960 2854.980 167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 215.960 2854.980 217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 265.960 2854.980 267.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 315.960 2854.980 317.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 365.960 2854.980 367.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 415.960 2854.980 417.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 465.960 2854.980 467.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 515.960 2854.980 517.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 565.960 2854.980 567.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 615.960 2854.980 617.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 665.960 2854.980 667.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 715.960 2854.980 717.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 765.960 2854.980 767.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 815.960 2854.980 817.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 865.960 2854.980 867.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 915.960 2854.980 917.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 965.960 2854.980 967.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1015.960 2854.980 1017.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1065.960 2854.980 1067.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1115.960 2854.980 1117.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1165.960 2854.980 1167.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1215.960 2854.980 1217.560 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1265.960 2854.980 1267.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.120 11.460 347.720 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 525.880 11.460 527.480 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 702.280 11.460 703.880 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 882.040 11.460 883.640 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1238.760 11.460 1240.360 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1596.040 11.460 1597.640 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1775.240 11.460 1776.840 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1952.760 11.460 1954.360 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2131.400 11.460 2133.000 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2488.680 11.460 2490.280 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2842.040 11.460 2843.640 1286.060 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 1.580 0.260 3.580 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 0.260 2854.980 2.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1307.020 2854.980 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2852.980 0.260 2854.980 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 0.260 19.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 17.580 1286.000 19.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.580 0.260 69.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 0.260 119.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.580 1286.000 119.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.580 0.260 169.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.580 0.260 219.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.580 1286.000 219.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 267.580 0.260 269.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 317.580 0.260 319.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 317.580 1286.000 319.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 367.580 0.260 369.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 367.580 1286.625 369.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 417.580 0.260 419.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 467.580 0.260 469.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 467.580 1286.625 469.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 517.580 0.260 519.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 567.580 0.260 569.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 617.580 0.260 619.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 617.580 1286.625 619.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 667.580 0.260 669.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 717.580 0.260 719.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 767.580 0.260 769.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 767.580 1286.000 769.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 817.580 0.260 819.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.580 0.260 869.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 917.580 0.260 919.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 967.580 0.260 969.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 967.580 1286.000 969.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1017.580 0.260 1019.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1067.580 0.260 1069.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1117.580 0.260 1119.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1117.580 1286.625 1119.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1167.580 0.260 1169.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1217.580 0.260 1219.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1217.580 1286.625 1219.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1267.580 0.260 1269.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1267.580 1286.625 1269.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1317.580 0.260 1319.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1367.580 0.260 1369.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1417.580 0.260 1419.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1467.580 0.260 1469.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1517.580 0.260 1519.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1517.580 1286.000 1519.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1567.580 0.260 1569.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1617.580 0.260 1619.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1617.580 1286.625 1619.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1667.580 0.260 1669.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1717.580 0.260 1719.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1717.580 1286.000 1719.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1767.580 0.260 1769.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1817.580 0.260 1819.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1867.580 0.260 1869.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1867.580 1286.000 1869.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1917.580 0.260 1919.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1967.580 0.260 1969.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2017.580 0.260 2019.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2067.580 0.260 2069.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2067.580 1286.000 2069.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2117.580 0.260 2119.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2167.580 0.260 2169.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2167.580 1286.000 2169.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2217.580 0.260 2219.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2217.580 1286.625 2219.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2267.580 0.260 2269.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2317.580 0.260 2319.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2367.580 0.260 2369.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2367.580 1286.000 2369.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2417.580 0.260 2419.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2467.580 0.260 2469.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2467.580 1286.625 2469.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2517.580 0.260 2519.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2517.580 1286.000 2519.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2567.580 0.260 2569.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2617.580 0.260 2619.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2617.580 1286.000 2619.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2667.580 0.260 2669.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2717.580 0.260 2719.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2717.580 1286.000 2719.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2767.580 0.260 2769.180 1309.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2817.580 0.260 2819.180 4.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2817.580 1286.000 2819.180 1309.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 19.260 2854.980 20.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 69.260 2854.980 70.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 119.260 2854.980 120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 169.260 2854.980 170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 219.260 2854.980 220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 269.260 2854.980 270.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 319.260 2854.980 320.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 369.260 2854.980 370.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 419.260 2854.980 420.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 469.260 2854.980 470.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 519.260 2854.980 520.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 569.260 2854.980 570.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 619.260 2854.980 620.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 669.260 2854.980 670.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 719.260 2854.980 720.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 769.260 2854.980 770.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 819.260 2854.980 820.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 869.260 2854.980 870.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 919.260 2854.980 920.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 969.260 2854.980 970.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1019.260 2854.980 1020.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1069.260 2854.980 1070.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1119.260 2854.980 1120.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1169.260 2854.980 1170.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1219.260 2854.980 1220.860 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1.580 1269.260 2854.980 1270.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 349.480 11.460 351.080 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 529.240 11.460 530.840 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 705.640 11.460 707.240 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 885.400 11.460 887.000 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1242.120 11.460 1243.720 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1599.400 11.460 1601.000 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1778.600 11.460 1780.200 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1956.120 11.460 1957.720 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2134.760 11.460 2136.360 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2492.040 11.460 2493.640 1286.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2844.280 11.460 2845.880 1286.060 ;
    END
  END VSS
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1310.505 84.560 1311.065 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 1310.505 218.960 1311.065 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 1310.505 252.560 1311.065 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1310.505 286.160 1311.065 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1310.505 319.760 1311.065 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 1310.505 353.360 1311.065 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1310.505 386.960 1311.065 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1310.505 420.560 1311.065 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1310.505 454.160 1311.065 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.816000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1310.505 487.760 1311.065 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1310.505 521.360 1311.065 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1310.505 151.760 1311.065 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1310.505 50.960 1311.065 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1310.505 554.960 1311.065 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 1310.505 890.960 1311.065 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 1310.505 924.560 1311.065 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 1310.505 958.160 1311.065 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 1310.505 991.760 1311.065 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1024.800 1310.505 1025.360 1311.065 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 1310.505 1058.960 1311.065 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 1310.505 1092.560 1311.065 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 1310.505 1126.160 1311.065 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 1310.505 1159.760 1311.065 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 1310.505 1193.360 1311.065 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 1310.505 588.560 1311.065 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1226.400 1310.505 1226.960 1311.065 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1260.000 1310.505 1260.560 1311.065 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1293.600 1310.505 1294.160 1311.065 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1327.200 1310.505 1327.760 1311.065 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1360.800 1310.505 1361.360 1311.065 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 1310.505 1394.960 1311.065 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1428.000 1310.505 1428.560 1311.065 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1461.600 1310.505 1462.160 1311.065 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1495.200 1310.505 1495.760 1311.065 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 1310.505 1529.360 1311.065 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1310.505 622.160 1311.065 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1562.400 1310.505 1562.960 1311.065 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1596.000 1310.505 1596.560 1311.065 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1310.505 655.760 1311.065 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 1310.505 689.360 1311.065 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 1310.505 722.960 1311.065 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 1310.505 756.560 1311.065 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1310.505 790.160 1311.065 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 1310.505 823.760 1311.065 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1310.505 857.360 1311.065 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 1310.505 1764.560 1311.065 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 1310.505 2100.560 1311.065 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2133.600 1310.505 2134.160 1311.065 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2167.200 1310.505 2167.760 1311.065 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2200.800 1310.505 2201.360 1311.065 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2234.400 1310.505 2234.960 1311.065 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2268.000 1310.505 2268.560 1311.065 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2301.600 1310.505 2302.160 1311.065 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2335.200 1310.505 2335.760 1311.065 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2368.800 1310.505 2369.360 1311.065 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2402.400 1310.505 2402.960 1311.065 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1797.600 1310.505 1798.160 1311.065 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2436.000 1310.505 2436.560 1311.065 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2469.600 1310.505 2470.160 1311.065 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2503.200 1310.505 2503.760 1311.065 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2536.800 1310.505 2537.360 1311.065 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2570.400 1310.505 2570.960 1311.065 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2604.000 1310.505 2604.560 1311.065 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2637.600 1310.505 2638.160 1311.065 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2671.200 1310.505 2671.760 1311.065 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2704.800 1310.505 2705.360 1311.065 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2738.400 1310.505 2738.960 1311.065 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1831.200 1310.505 1831.760 1311.065 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2772.000 1310.505 2772.560 1311.065 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2805.600 1310.505 2806.160 1311.065 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1864.800 1310.505 1865.360 1311.065 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1898.400 1310.505 1898.960 1311.065 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1932.000 1310.505 1932.560 1311.065 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1965.600 1310.505 1966.160 1311.065 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 1999.200 1310.505 1999.760 1311.065 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2032.800 1310.505 2033.360 1311.065 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal2 ;
        RECT 2066.400 1310.505 2066.960 1311.065 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 1310.505 118.160 1311.065 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 1310.505 1630.160 1311.065 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 1310.505 1663.760 1311.065 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 1310.505 1697.360 1311.065 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1730.400 1310.505 1730.960 1311.065 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1310.505 17.360 1311.065 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1310.505 185.360 1311.065 ;
    END
  END wb_we_i
  PIN write_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1128.447998 ;
    ANTENNADIFFAREA 210.124802 ;
    PORT
      LAYER Metal2 ;
        RECT 2839.200 1310.505 2839.760 1311.065 ;
    END
  END write_enable_i
  OBS
      LAYER Nwell ;
        RECT 9.650 11.330 2846.910 1297.950 ;
      LAYER Metal1 ;
        RECT 10.080 11.460 2846.480 1297.820 ;
      LAYER Metal2 ;
        RECT 9.100 1310.205 16.500 1310.820 ;
        RECT 17.660 1310.205 50.100 1310.820 ;
        RECT 51.260 1310.205 83.700 1310.820 ;
        RECT 84.860 1310.205 117.300 1310.820 ;
        RECT 118.460 1310.205 150.900 1310.820 ;
        RECT 152.060 1310.205 184.500 1310.820 ;
        RECT 185.660 1310.205 218.100 1310.820 ;
        RECT 219.260 1310.205 251.700 1310.820 ;
        RECT 252.860 1310.205 285.300 1310.820 ;
        RECT 286.460 1310.205 318.900 1310.820 ;
        RECT 320.060 1310.205 352.500 1310.820 ;
        RECT 353.660 1310.205 386.100 1310.820 ;
        RECT 387.260 1310.205 419.700 1310.820 ;
        RECT 420.860 1310.205 453.300 1310.820 ;
        RECT 454.460 1310.205 486.900 1310.820 ;
        RECT 488.060 1310.205 520.500 1310.820 ;
        RECT 521.660 1310.205 554.100 1310.820 ;
        RECT 555.260 1310.205 587.700 1310.820 ;
        RECT 588.860 1310.205 621.300 1310.820 ;
        RECT 622.460 1310.205 654.900 1310.820 ;
        RECT 656.060 1310.205 688.500 1310.820 ;
        RECT 689.660 1310.205 722.100 1310.820 ;
        RECT 723.260 1310.205 755.700 1310.820 ;
        RECT 756.860 1310.205 789.300 1310.820 ;
        RECT 790.460 1310.205 822.900 1310.820 ;
        RECT 824.060 1310.205 856.500 1310.820 ;
        RECT 857.660 1310.205 890.100 1310.820 ;
        RECT 891.260 1310.205 923.700 1310.820 ;
        RECT 924.860 1310.205 957.300 1310.820 ;
        RECT 958.460 1310.205 990.900 1310.820 ;
        RECT 992.060 1310.205 1024.500 1310.820 ;
        RECT 1025.660 1310.205 1058.100 1310.820 ;
        RECT 1059.260 1310.205 1091.700 1310.820 ;
        RECT 1092.860 1310.205 1125.300 1310.820 ;
        RECT 1126.460 1310.205 1158.900 1310.820 ;
        RECT 1160.060 1310.205 1192.500 1310.820 ;
        RECT 1193.660 1310.205 1226.100 1310.820 ;
        RECT 1227.260 1310.205 1259.700 1310.820 ;
        RECT 1260.860 1310.205 1293.300 1310.820 ;
        RECT 1294.460 1310.205 1326.900 1310.820 ;
        RECT 1328.060 1310.205 1360.500 1310.820 ;
        RECT 1361.660 1310.205 1394.100 1310.820 ;
        RECT 1395.260 1310.205 1427.700 1310.820 ;
        RECT 1428.860 1310.205 1461.300 1310.820 ;
        RECT 1462.460 1310.205 1494.900 1310.820 ;
        RECT 1496.060 1310.205 1528.500 1310.820 ;
        RECT 1529.660 1310.205 1562.100 1310.820 ;
        RECT 1563.260 1310.205 1595.700 1310.820 ;
        RECT 1596.860 1310.205 1629.300 1310.820 ;
        RECT 1630.460 1310.205 1662.900 1310.820 ;
        RECT 1664.060 1310.205 1696.500 1310.820 ;
        RECT 1697.660 1310.205 1730.100 1310.820 ;
        RECT 1731.260 1310.205 1763.700 1310.820 ;
        RECT 1764.860 1310.205 1797.300 1310.820 ;
        RECT 1798.460 1310.205 1830.900 1310.820 ;
        RECT 1832.060 1310.205 1864.500 1310.820 ;
        RECT 1865.660 1310.205 1898.100 1310.820 ;
        RECT 1899.260 1310.205 1931.700 1310.820 ;
        RECT 1932.860 1310.205 1965.300 1310.820 ;
        RECT 1966.460 1310.205 1998.900 1310.820 ;
        RECT 2000.060 1310.205 2032.500 1310.820 ;
        RECT 2033.660 1310.205 2066.100 1310.820 ;
        RECT 2067.260 1310.205 2099.700 1310.820 ;
        RECT 2100.860 1310.205 2133.300 1310.820 ;
        RECT 2134.460 1310.205 2166.900 1310.820 ;
        RECT 2168.060 1310.205 2200.500 1310.820 ;
        RECT 2201.660 1310.205 2234.100 1310.820 ;
        RECT 2235.260 1310.205 2267.700 1310.820 ;
        RECT 2268.860 1310.205 2301.300 1310.820 ;
        RECT 2302.460 1310.205 2334.900 1310.820 ;
        RECT 2336.060 1310.205 2368.500 1310.820 ;
        RECT 2369.660 1310.205 2402.100 1310.820 ;
        RECT 2403.260 1310.205 2435.700 1310.820 ;
        RECT 2436.860 1310.205 2469.300 1310.820 ;
        RECT 2470.460 1310.205 2502.900 1310.820 ;
        RECT 2504.060 1310.205 2536.500 1310.820 ;
        RECT 2537.660 1310.205 2570.100 1310.820 ;
        RECT 2571.260 1310.205 2603.700 1310.820 ;
        RECT 2604.860 1310.205 2637.300 1310.820 ;
        RECT 2638.460 1310.205 2670.900 1310.820 ;
        RECT 2672.060 1310.205 2704.500 1310.820 ;
        RECT 2705.660 1310.205 2738.100 1310.820 ;
        RECT 2739.260 1310.205 2771.700 1310.820 ;
        RECT 2772.860 1310.205 2805.300 1310.820 ;
        RECT 2806.460 1310.205 2838.900 1310.820 ;
        RECT 2840.060 1310.205 2845.740 1310.820 ;
        RECT 9.100 1.210 2845.740 1310.205 ;
      LAYER Metal3 ;
        RECT 9.050 1.260 2845.790 1309.700 ;
      LAYER Metal4 ;
        RECT 10.240 1286.325 13.980 1309.190 ;
        RECT 16.180 1286.325 17.280 1309.190 ;
        RECT 10.240 1285.700 17.280 1286.325 ;
        RECT 19.480 1285.700 63.980 1309.190 ;
        RECT 10.240 4.740 63.980 1285.700 ;
        RECT 10.240 1.210 13.980 4.740 ;
        RECT 16.180 1.210 17.280 4.740 ;
        RECT 19.480 1.210 63.980 4.740 ;
        RECT 66.180 1.210 67.280 1309.190 ;
        RECT 69.480 1285.280 113.980 1309.190 ;
        RECT 116.180 1285.700 117.280 1309.190 ;
        RECT 119.480 1285.700 163.980 1309.190 ;
        RECT 116.180 1285.280 163.980 1285.700 ;
        RECT 69.480 4.740 163.980 1285.280 ;
        RECT 69.480 1.210 113.980 4.740 ;
        RECT 116.180 1.210 117.280 4.740 ;
        RECT 119.480 1.210 163.980 4.740 ;
        RECT 166.180 1.210 167.280 1309.190 ;
        RECT 169.480 1.210 213.980 1309.190 ;
        RECT 216.180 1285.700 217.280 1309.190 ;
        RECT 219.480 1285.700 263.980 1309.190 ;
        RECT 216.180 4.740 263.980 1285.700 ;
        RECT 216.180 1.210 217.280 4.740 ;
        RECT 219.480 1.210 263.980 4.740 ;
        RECT 266.180 1.210 267.280 1309.190 ;
        RECT 269.480 1285.280 313.980 1309.190 ;
        RECT 316.180 1285.700 317.280 1309.190 ;
        RECT 319.480 1286.360 363.980 1309.190 ;
        RECT 319.480 1285.700 345.820 1286.360 ;
        RECT 316.180 1285.280 345.820 1285.700 ;
        RECT 269.480 11.160 345.820 1285.280 ;
        RECT 348.020 11.160 349.180 1286.360 ;
        RECT 351.380 11.160 363.980 1286.360 ;
        RECT 269.480 4.740 363.980 11.160 ;
        RECT 269.480 1.210 313.980 4.740 ;
        RECT 316.180 1.210 317.280 4.740 ;
        RECT 319.480 1.210 363.980 4.740 ;
        RECT 366.180 1286.325 367.280 1309.190 ;
        RECT 369.480 1286.325 413.980 1309.190 ;
        RECT 366.180 1285.280 413.980 1286.325 ;
        RECT 416.180 1285.280 417.280 1309.190 ;
        RECT 366.180 4.740 417.280 1285.280 ;
        RECT 366.180 1.210 367.280 4.740 ;
        RECT 369.480 1.210 413.980 4.740 ;
        RECT 416.180 1.210 417.280 4.740 ;
        RECT 419.480 1.210 463.980 1309.190 ;
        RECT 466.180 1286.325 467.280 1309.190 ;
        RECT 469.480 1286.325 513.980 1309.190 ;
        RECT 466.180 4.740 513.980 1286.325 ;
        RECT 466.180 1.210 467.280 4.740 ;
        RECT 469.480 1.210 513.980 4.740 ;
        RECT 516.180 1.210 517.280 1309.190 ;
        RECT 519.480 1286.360 563.980 1309.190 ;
        RECT 519.480 11.160 525.580 1286.360 ;
        RECT 527.780 11.160 528.940 1286.360 ;
        RECT 531.140 11.160 563.980 1286.360 ;
        RECT 519.480 1.210 563.980 11.160 ;
        RECT 566.180 1.210 567.280 1309.190 ;
        RECT 569.480 1285.280 613.980 1309.190 ;
        RECT 616.180 1286.325 617.280 1309.190 ;
        RECT 619.480 1286.325 663.980 1309.190 ;
        RECT 616.180 1285.280 663.980 1286.325 ;
        RECT 569.480 4.740 663.980 1285.280 ;
        RECT 569.480 1.210 613.980 4.740 ;
        RECT 616.180 1.210 617.280 4.740 ;
        RECT 619.480 1.210 663.980 4.740 ;
        RECT 666.180 1.210 667.280 1309.190 ;
        RECT 669.480 1286.360 713.980 1309.190 ;
        RECT 669.480 11.160 701.980 1286.360 ;
        RECT 704.180 11.160 705.340 1286.360 ;
        RECT 707.540 11.160 713.980 1286.360 ;
        RECT 669.480 1.210 713.980 11.160 ;
        RECT 716.180 1.210 717.280 1309.190 ;
        RECT 719.480 1285.280 763.980 1309.190 ;
        RECT 766.180 1285.700 767.280 1309.190 ;
        RECT 769.480 1285.700 813.980 1309.190 ;
        RECT 766.180 1285.280 813.980 1285.700 ;
        RECT 719.480 4.740 813.980 1285.280 ;
        RECT 719.480 1.210 763.980 4.740 ;
        RECT 766.180 1.210 767.280 4.740 ;
        RECT 769.480 1.210 813.980 4.740 ;
        RECT 816.180 1.210 817.280 1309.190 ;
        RECT 819.480 1286.325 863.980 1309.190 ;
        RECT 866.180 1286.325 867.280 1309.190 ;
        RECT 819.480 4.740 867.280 1286.325 ;
        RECT 819.480 1.210 863.980 4.740 ;
        RECT 866.180 1.210 867.280 4.740 ;
        RECT 869.480 1286.360 913.980 1309.190 ;
        RECT 869.480 11.160 881.740 1286.360 ;
        RECT 883.940 11.160 885.100 1286.360 ;
        RECT 887.300 11.160 913.980 1286.360 ;
        RECT 869.480 1.210 913.980 11.160 ;
        RECT 916.180 1.210 917.280 1309.190 ;
        RECT 919.480 1285.280 963.980 1309.190 ;
        RECT 966.180 1285.700 967.280 1309.190 ;
        RECT 969.480 1285.700 1013.980 1309.190 ;
        RECT 966.180 1285.280 1013.980 1285.700 ;
        RECT 919.480 4.740 1013.980 1285.280 ;
        RECT 919.480 1.210 963.980 4.740 ;
        RECT 966.180 1.210 967.280 4.740 ;
        RECT 969.480 1.210 1013.980 4.740 ;
        RECT 1016.180 1.210 1017.280 1309.190 ;
        RECT 1019.480 1.210 1063.980 1309.190 ;
        RECT 1066.180 1.210 1067.280 1309.190 ;
        RECT 1069.480 1286.325 1113.980 1309.190 ;
        RECT 1116.180 1286.325 1117.280 1309.190 ;
        RECT 1119.480 1286.325 1163.980 1309.190 ;
        RECT 1069.480 4.740 1163.980 1286.325 ;
        RECT 1069.480 1.210 1113.980 4.740 ;
        RECT 1116.180 1.210 1117.280 4.740 ;
        RECT 1119.480 1.210 1163.980 4.740 ;
        RECT 1166.180 1.210 1167.280 1309.190 ;
        RECT 1169.480 1286.325 1213.980 1309.190 ;
        RECT 1216.180 1286.325 1217.280 1309.190 ;
        RECT 1219.480 1286.360 1263.980 1309.190 ;
        RECT 1219.480 1286.325 1238.460 1286.360 ;
        RECT 1169.480 11.160 1238.460 1286.325 ;
        RECT 1240.660 11.160 1241.820 1286.360 ;
        RECT 1244.020 1286.325 1263.980 1286.360 ;
        RECT 1266.180 1286.325 1267.280 1309.190 ;
        RECT 1269.480 1286.325 1313.980 1309.190 ;
        RECT 1244.020 11.160 1313.980 1286.325 ;
        RECT 1169.480 4.740 1313.980 11.160 ;
        RECT 1169.480 1.210 1213.980 4.740 ;
        RECT 1216.180 1.210 1217.280 4.740 ;
        RECT 1219.480 1.210 1263.980 4.740 ;
        RECT 1266.180 1.210 1267.280 4.740 ;
        RECT 1269.480 1.210 1313.980 4.740 ;
        RECT 1316.180 1.210 1317.280 1309.190 ;
        RECT 1319.480 1286.325 1363.980 1309.190 ;
        RECT 1366.180 1286.325 1367.280 1309.190 ;
        RECT 1319.480 4.740 1367.280 1286.325 ;
        RECT 1319.480 1.210 1363.980 4.740 ;
        RECT 1366.180 1.210 1367.280 4.740 ;
        RECT 1369.480 1.210 1413.980 1309.190 ;
        RECT 1416.180 1.210 1417.280 1309.190 ;
        RECT 1419.480 1.210 1463.980 1309.190 ;
        RECT 1466.180 1.210 1467.280 1309.190 ;
        RECT 1469.480 1285.280 1513.980 1309.190 ;
        RECT 1516.180 1285.700 1517.280 1309.190 ;
        RECT 1519.480 1285.700 1563.980 1309.190 ;
        RECT 1516.180 1285.280 1563.980 1285.700 ;
        RECT 1469.480 4.740 1563.980 1285.280 ;
        RECT 1469.480 1.210 1513.980 4.740 ;
        RECT 1516.180 1.210 1517.280 4.740 ;
        RECT 1519.480 1.210 1563.980 4.740 ;
        RECT 1566.180 1.210 1567.280 1309.190 ;
        RECT 1569.480 1286.360 1613.980 1309.190 ;
        RECT 1569.480 11.160 1595.740 1286.360 ;
        RECT 1597.940 11.160 1599.100 1286.360 ;
        RECT 1601.300 11.160 1613.980 1286.360 ;
        RECT 1569.480 1.210 1613.980 11.160 ;
        RECT 1616.180 1286.325 1617.280 1309.190 ;
        RECT 1619.480 1286.325 1663.980 1309.190 ;
        RECT 1616.180 4.740 1663.980 1286.325 ;
        RECT 1616.180 1.210 1617.280 4.740 ;
        RECT 1619.480 1.210 1663.980 4.740 ;
        RECT 1666.180 1.210 1667.280 1309.190 ;
        RECT 1669.480 1285.280 1713.980 1309.190 ;
        RECT 1716.180 1285.700 1717.280 1309.190 ;
        RECT 1719.480 1285.700 1763.980 1309.190 ;
        RECT 1716.180 1285.280 1763.980 1285.700 ;
        RECT 1669.480 4.740 1763.980 1285.280 ;
        RECT 1669.480 1.210 1713.980 4.740 ;
        RECT 1716.180 1.210 1717.280 4.740 ;
        RECT 1719.480 1.210 1763.980 4.740 ;
        RECT 1766.180 1.210 1767.280 1309.190 ;
        RECT 1769.480 1286.360 1813.980 1309.190 ;
        RECT 1769.480 11.160 1774.940 1286.360 ;
        RECT 1777.140 11.160 1778.300 1286.360 ;
        RECT 1780.500 11.160 1813.980 1286.360 ;
        RECT 1769.480 1.210 1813.980 11.160 ;
        RECT 1816.180 1.210 1817.280 1309.190 ;
        RECT 1819.480 1286.325 1863.980 1309.190 ;
        RECT 1866.180 1286.325 1867.280 1309.190 ;
        RECT 1819.480 1285.700 1867.280 1286.325 ;
        RECT 1869.480 1285.700 1913.980 1309.190 ;
        RECT 1819.480 4.740 1913.980 1285.700 ;
        RECT 1819.480 1.210 1863.980 4.740 ;
        RECT 1866.180 1.210 1867.280 4.740 ;
        RECT 1869.480 1.210 1913.980 4.740 ;
        RECT 1916.180 1.210 1917.280 1309.190 ;
        RECT 1919.480 1286.360 1963.980 1309.190 ;
        RECT 1919.480 11.160 1952.460 1286.360 ;
        RECT 1954.660 11.160 1955.820 1286.360 ;
        RECT 1958.020 11.160 1963.980 1286.360 ;
        RECT 1919.480 1.210 1963.980 11.160 ;
        RECT 1966.180 1.210 1967.280 1309.190 ;
        RECT 1969.480 1286.325 2013.980 1309.190 ;
        RECT 2016.180 1286.325 2017.280 1309.190 ;
        RECT 1969.480 4.740 2017.280 1286.325 ;
        RECT 1969.480 1.210 2013.980 4.740 ;
        RECT 2016.180 1.210 2017.280 4.740 ;
        RECT 2019.480 1.210 2063.980 1309.190 ;
        RECT 2066.180 1285.700 2067.280 1309.190 ;
        RECT 2069.480 1286.325 2113.980 1309.190 ;
        RECT 2116.180 1286.325 2117.280 1309.190 ;
        RECT 2069.480 1285.700 2117.280 1286.325 ;
        RECT 2066.180 4.740 2117.280 1285.700 ;
        RECT 2066.180 1.210 2067.280 4.740 ;
        RECT 2069.480 1.210 2113.980 4.740 ;
        RECT 2116.180 1.210 2117.280 4.740 ;
        RECT 2119.480 1286.360 2163.980 1309.190 ;
        RECT 2119.480 11.160 2131.100 1286.360 ;
        RECT 2133.300 11.160 2134.460 1286.360 ;
        RECT 2136.660 1285.280 2163.980 1286.360 ;
        RECT 2166.180 1285.700 2167.280 1309.190 ;
        RECT 2169.480 1285.700 2213.980 1309.190 ;
        RECT 2166.180 1285.280 2213.980 1285.700 ;
        RECT 2136.660 11.160 2213.980 1285.280 ;
        RECT 2119.480 4.740 2213.980 11.160 ;
        RECT 2119.480 1.210 2163.980 4.740 ;
        RECT 2166.180 1.210 2167.280 4.740 ;
        RECT 2169.480 1.210 2213.980 4.740 ;
        RECT 2216.180 1286.325 2217.280 1309.190 ;
        RECT 2219.480 1286.325 2263.980 1309.190 ;
        RECT 2216.180 1285.280 2263.980 1286.325 ;
        RECT 2266.180 1285.280 2267.280 1309.190 ;
        RECT 2216.180 4.740 2267.280 1285.280 ;
        RECT 2216.180 1.210 2217.280 4.740 ;
        RECT 2219.480 1.210 2263.980 4.740 ;
        RECT 2266.180 1.210 2267.280 4.740 ;
        RECT 2269.480 1.210 2313.980 1309.190 ;
        RECT 2316.180 1.210 2317.280 1309.190 ;
        RECT 2319.480 1285.280 2363.980 1309.190 ;
        RECT 2366.180 1285.700 2367.280 1309.190 ;
        RECT 2369.480 1285.700 2413.980 1309.190 ;
        RECT 2366.180 1285.280 2413.980 1285.700 ;
        RECT 2319.480 4.740 2413.980 1285.280 ;
        RECT 2319.480 1.210 2363.980 4.740 ;
        RECT 2366.180 1.210 2367.280 4.740 ;
        RECT 2369.480 1.210 2413.980 4.740 ;
        RECT 2416.180 1.210 2417.280 1309.190 ;
        RECT 2419.480 1285.280 2463.980 1309.190 ;
        RECT 2466.180 1286.325 2467.280 1309.190 ;
        RECT 2469.480 1286.360 2513.980 1309.190 ;
        RECT 2469.480 1286.325 2488.380 1286.360 ;
        RECT 2466.180 1285.280 2488.380 1286.325 ;
        RECT 2419.480 11.160 2488.380 1285.280 ;
        RECT 2490.580 11.160 2491.740 1286.360 ;
        RECT 2493.940 1286.325 2513.980 1286.360 ;
        RECT 2516.180 1286.325 2517.280 1309.190 ;
        RECT 2493.940 1285.700 2517.280 1286.325 ;
        RECT 2519.480 1285.700 2563.980 1309.190 ;
        RECT 2493.940 11.160 2563.980 1285.700 ;
        RECT 2419.480 4.740 2563.980 11.160 ;
        RECT 2419.480 1.210 2463.980 4.740 ;
        RECT 2466.180 1.210 2467.280 4.740 ;
        RECT 2469.480 1.210 2513.980 4.740 ;
        RECT 2516.180 1.210 2517.280 4.740 ;
        RECT 2519.480 1.210 2563.980 4.740 ;
        RECT 2566.180 1.210 2567.280 1309.190 ;
        RECT 2569.480 1285.280 2613.980 1309.190 ;
        RECT 2616.180 1285.700 2617.280 1309.190 ;
        RECT 2619.480 1285.700 2663.980 1309.190 ;
        RECT 2616.180 1285.280 2663.980 1285.700 ;
        RECT 2569.480 4.740 2663.980 1285.280 ;
        RECT 2569.480 1.210 2613.980 4.740 ;
        RECT 2616.180 1.210 2617.280 4.740 ;
        RECT 2619.480 1.210 2663.980 4.740 ;
        RECT 2666.180 1.210 2667.280 1309.190 ;
        RECT 2669.480 1285.280 2713.980 1309.190 ;
        RECT 2716.180 1285.700 2717.280 1309.190 ;
        RECT 2719.480 1285.700 2763.980 1309.190 ;
        RECT 2716.180 1285.280 2763.980 1285.700 ;
        RECT 2669.480 4.740 2763.980 1285.280 ;
        RECT 2669.480 1.210 2713.980 4.740 ;
        RECT 2716.180 1.210 2717.280 4.740 ;
        RECT 2719.480 1.210 2763.980 4.740 ;
        RECT 2766.180 1.210 2767.280 1309.190 ;
        RECT 2769.480 1285.280 2813.980 1309.190 ;
        RECT 2816.180 1285.700 2817.280 1309.190 ;
        RECT 2819.480 1285.700 2839.060 1309.190 ;
        RECT 2816.180 1285.280 2839.060 1285.700 ;
        RECT 2769.480 4.740 2839.060 1285.280 ;
        RECT 2769.480 1.210 2813.980 4.740 ;
        RECT 2816.180 1.210 2817.280 4.740 ;
        RECT 2819.480 1.210 2839.060 4.740 ;
  END
END efuse_wb_mem_1024x32
END LIBRARY

