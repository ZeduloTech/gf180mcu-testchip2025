VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2900.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 14.080 17.440 24.080 982.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 17.440 2884.480 27.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 972.160 2884.480 982.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2874.480 17.440 2884.480 982.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.080 5.440 29.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.080 5.440 109.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.080 5.440 189.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.080 5.440 269.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.080 5.440 349.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.080 5.440 429.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.080 5.440 509.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.080 5.440 589.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 5.440 669.080 66.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 545.800 669.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.080 5.440 749.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.080 5.440 829.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.080 5.440 909.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 5.440 989.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.080 5.440 1069.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.080 5.440 1149.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.080 5.440 1229.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.080 5.440 1309.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.080 5.440 1389.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.080 5.440 1469.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 5.440 1549.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.080 5.440 1629.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.080 5.440 1709.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.080 5.440 1789.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.080 5.440 1869.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.080 5.440 1949.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.080 5.440 2029.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.080 5.440 2109.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.080 5.440 2189.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.080 5.440 2269.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.080 5.440 2349.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 5.440 2429.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 5.440 2509.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 5.440 2589.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 5.440 2669.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 144.725 2669.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 5.440 2749.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 5.440 2829.080 994.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 56.590 2896.480 59.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 116.590 2635.895 119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 176.590 2896.480 179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 236.590 2896.480 239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 296.590 2896.480 299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 356.590 2896.480 359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 416.590 2896.480 419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 476.590 2896.480 479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 536.590 2896.480 539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 596.590 2896.480 599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 656.590 2896.480 659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 716.590 2896.480 719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 776.590 2896.480 779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 836.590 2896.480 839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 896.590 2896.480 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 956.590 2896.480 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 116.590 2896.480 119.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2620.580 5.440 2623.580 994.160 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 2.080 5.440 12.080 994.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 5.440 2896.480 15.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 984.160 2896.480 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2886.480 5.440 2896.480 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 48.080 5.440 51.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 5.440 131.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.080 5.440 211.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.080 5.440 291.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.080 5.440 371.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.080 5.440 451.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 528.080 5.440 531.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 608.080 5.440 611.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.080 5.440 691.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 768.080 5.440 771.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 848.080 5.440 851.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.080 5.440 931.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1008.080 5.440 1011.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 5.440 1091.080 66.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 545.800 1091.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1168.080 5.440 1171.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.080 5.440 1251.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1328.080 5.440 1331.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1408.080 5.440 1411.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1488.080 5.440 1491.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.080 5.440 1571.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.080 5.440 1651.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1728.080 5.440 1731.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1808.080 5.440 1811.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1888.080 5.440 1891.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.080 5.440 1971.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2048.080 5.440 2051.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2128.080 5.440 2131.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2208.080 5.440 2211.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2288.080 5.440 2291.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.080 5.440 2371.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 5.440 2451.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 5.440 2531.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 5.440 2611.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 5.440 2691.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 144.725 2691.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 5.440 2771.080 994.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 5.440 2851.080 994.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 86.590 2636.395 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 146.590 2635.895 149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 206.590 2896.480 209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 266.590 2896.480 269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 326.590 2896.480 329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 386.590 2896.480 389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 446.590 2896.480 449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 506.590 2896.480 509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 566.590 2896.480 569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 626.590 2896.480 629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 686.590 2896.480 689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 746.590 2896.480 749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 806.590 2896.480 809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 866.590 2896.480 869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 926.590 2896.480 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 86.590 2896.480 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 146.590 2896.480 149.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2632.580 5.440 2635.580 994.160 ;
    END
  END VSS
  PIN caravel_io_ie[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 0.560 ;
    END
  END caravel_io_ie[0]
  PIN caravel_io_ie[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 2242.240 0.000 2242.800 0.560 ;
    END
  END caravel_io_ie[10]
  PIN caravel_io_ie[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2457.280 0.000 2457.840 0.560 ;
    END
  END caravel_io_ie[11]
  PIN caravel_io_ie[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2672.320 0.000 2672.880 0.560 ;
    END
  END caravel_io_ie[12]
  PIN caravel_io_ie[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 0.560 ;
    END
  END caravel_io_ie[1]
  PIN caravel_io_ie[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 0.560 ;
    END
  END caravel_io_ie[2]
  PIN caravel_io_ie[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 0.000 737.520 0.560 ;
    END
  END caravel_io_ie[3]
  PIN caravel_io_ie[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 0.000 952.560 0.560 ;
    END
  END caravel_io_ie[4]
  PIN caravel_io_ie[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1167.040 0.000 1167.600 0.560 ;
    END
  END caravel_io_ie[5]
  PIN caravel_io_ie[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1382.080 0.000 1382.640 0.560 ;
    END
  END caravel_io_ie[6]
  PIN caravel_io_ie[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1597.120 0.000 1597.680 0.560 ;
    END
  END caravel_io_ie[7]
  PIN caravel_io_ie[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1812.160 0.000 1812.720 0.560 ;
    END
  END caravel_io_ie[8]
  PIN caravel_io_ie[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2027.200 0.000 2027.760 0.560 ;
    END
  END caravel_io_ie[9]
  PIN caravel_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 0.560 ;
    END
  END caravel_io_in[0]
  PIN caravel_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.867500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2269.120 0.000 2269.680 0.560 ;
    END
  END caravel_io_in[10]
  PIN caravel_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    PORT
      LAYER Metal2 ;
        RECT 2484.160 0.000 2484.720 0.560 ;
    END
  END caravel_io_in[11]
  PIN caravel_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2699.200 0.000 2699.760 0.560 ;
    END
  END caravel_io_in[12]
  PIN caravel_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 0.560 ;
    END
  END caravel_io_in[1]
  PIN caravel_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 0.560 ;
    END
  END caravel_io_in[2]
  PIN caravel_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 0.560 ;
    END
  END caravel_io_in[3]
  PIN caravel_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 978.880 0.000 979.440 0.560 ;
    END
  END caravel_io_in[4]
  PIN caravel_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 1193.920 0.000 1194.480 0.560 ;
    END
  END caravel_io_in[5]
  PIN caravel_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 1408.960 0.000 1409.520 0.560 ;
    END
  END caravel_io_in[6]
  PIN caravel_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 1624.000 0.000 1624.560 0.560 ;
    END
  END caravel_io_in[7]
  PIN caravel_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.867500 ;
    PORT
      LAYER Metal2 ;
        RECT 1839.040 0.000 1839.600 0.560 ;
    END
  END caravel_io_in[8]
  PIN caravel_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.867500 ;
    PORT
      LAYER Metal2 ;
        RECT 2054.080 0.000 2054.640 0.560 ;
    END
  END caravel_io_in[9]
  PIN caravel_io_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 0.560 ;
    END
  END caravel_io_oe[0]
  PIN caravel_io_oe[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2296.000 0.000 2296.560 0.560 ;
    END
  END caravel_io_oe[10]
  PIN caravel_io_oe[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2511.040 0.000 2511.600 0.560 ;
    END
  END caravel_io_oe[11]
  PIN caravel_io_oe[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2726.080 0.000 2726.640 0.560 ;
    END
  END caravel_io_oe[12]
  PIN caravel_io_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 0.560 ;
    END
  END caravel_io_oe[1]
  PIN caravel_io_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 0.560 ;
    END
  END caravel_io_oe[2]
  PIN caravel_io_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 0.560 ;
    END
  END caravel_io_oe[3]
  PIN caravel_io_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1005.760 0.000 1006.320 0.560 ;
    END
  END caravel_io_oe[4]
  PIN caravel_io_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1220.800 0.000 1221.360 0.560 ;
    END
  END caravel_io_oe[5]
  PIN caravel_io_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1435.840 0.000 1436.400 0.560 ;
    END
  END caravel_io_oe[6]
  PIN caravel_io_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1650.880 0.000 1651.440 0.560 ;
    END
  END caravel_io_oe[7]
  PIN caravel_io_oe[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1865.920 0.000 1866.480 0.560 ;
    END
  END caravel_io_oe[8]
  PIN caravel_io_oe[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2080.960 0.000 2081.520 0.560 ;
    END
  END caravel_io_oe[9]
  PIN caravel_io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 0.560 ;
    END
  END caravel_io_out[0]
  PIN caravel_io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2322.880 0.000 2323.440 0.560 ;
    END
  END caravel_io_out[10]
  PIN caravel_io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2537.920 0.000 2538.480 0.560 ;
    END
  END caravel_io_out[11]
  PIN caravel_io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2752.960 0.000 2753.520 0.560 ;
    END
  END caravel_io_out[12]
  PIN caravel_io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 0.560 ;
    END
  END caravel_io_out[1]
  PIN caravel_io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 0.560 ;
    END
  END caravel_io_out[2]
  PIN caravel_io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 0.560 ;
    END
  END caravel_io_out[3]
  PIN caravel_io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1032.640 0.000 1033.200 0.560 ;
    END
  END caravel_io_out[4]
  PIN caravel_io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1247.680 0.000 1248.240 0.560 ;
    END
  END caravel_io_out[5]
  PIN caravel_io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1462.720 0.000 1463.280 0.560 ;
    END
  END caravel_io_out[6]
  PIN caravel_io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1677.760 0.000 1678.320 0.560 ;
    END
  END caravel_io_out[7]
  PIN caravel_io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1892.800 0.000 1893.360 0.560 ;
    END
  END caravel_io_out[8]
  PIN caravel_io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2107.840 0.000 2108.400 0.560 ;
    END
  END caravel_io_out[9]
  PIN caravel_io_pulldown_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 0.560 ;
    END
  END caravel_io_pulldown_sel[0]
  PIN caravel_io_pulldown_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2349.760 0.000 2350.320 0.560 ;
    END
  END caravel_io_pulldown_sel[10]
  PIN caravel_io_pulldown_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2564.800 0.000 2565.360 0.560 ;
    END
  END caravel_io_pulldown_sel[11]
  PIN caravel_io_pulldown_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2779.840 0.000 2780.400 0.560 ;
    END
  END caravel_io_pulldown_sel[12]
  PIN caravel_io_pulldown_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 0.560 ;
    END
  END caravel_io_pulldown_sel[1]
  PIN caravel_io_pulldown_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 0.000 630.000 0.560 ;
    END
  END caravel_io_pulldown_sel[2]
  PIN caravel_io_pulldown_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 844.480 0.000 845.040 0.560 ;
    END
  END caravel_io_pulldown_sel[3]
  PIN caravel_io_pulldown_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1059.520 0.000 1060.080 0.560 ;
    END
  END caravel_io_pulldown_sel[4]
  PIN caravel_io_pulldown_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1274.560 0.000 1275.120 0.560 ;
    END
  END caravel_io_pulldown_sel[5]
  PIN caravel_io_pulldown_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1489.600 0.000 1490.160 0.560 ;
    END
  END caravel_io_pulldown_sel[6]
  PIN caravel_io_pulldown_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1704.640 0.000 1705.200 0.560 ;
    END
  END caravel_io_pulldown_sel[7]
  PIN caravel_io_pulldown_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1919.680 0.000 1920.240 0.560 ;
    END
  END caravel_io_pulldown_sel[8]
  PIN caravel_io_pulldown_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2134.720 0.000 2135.280 0.560 ;
    END
  END caravel_io_pulldown_sel[9]
  PIN caravel_io_pullup_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 0.560 ;
    END
  END caravel_io_pullup_sel[0]
  PIN caravel_io_pullup_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2376.640 0.000 2377.200 0.560 ;
    END
  END caravel_io_pullup_sel[10]
  PIN caravel_io_pullup_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2591.680 0.000 2592.240 0.560 ;
    END
  END caravel_io_pullup_sel[11]
  PIN caravel_io_pullup_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2806.720 0.000 2807.280 0.560 ;
    END
  END caravel_io_pullup_sel[12]
  PIN caravel_io_pullup_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 0.560 ;
    END
  END caravel_io_pullup_sel[1]
  PIN caravel_io_pullup_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 0.560 ;
    END
  END caravel_io_pullup_sel[2]
  PIN caravel_io_pullup_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 0.000 871.920 0.560 ;
    END
  END caravel_io_pullup_sel[3]
  PIN caravel_io_pullup_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1086.400 0.000 1086.960 0.560 ;
    END
  END caravel_io_pullup_sel[4]
  PIN caravel_io_pullup_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1301.440 0.000 1302.000 0.560 ;
    END
  END caravel_io_pullup_sel[5]
  PIN caravel_io_pullup_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1516.480 0.000 1517.040 0.560 ;
    END
  END caravel_io_pullup_sel[6]
  PIN caravel_io_pullup_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1731.520 0.000 1732.080 0.560 ;
    END
  END caravel_io_pullup_sel[7]
  PIN caravel_io_pullup_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1946.560 0.000 1947.120 0.560 ;
    END
  END caravel_io_pullup_sel[8]
  PIN caravel_io_pullup_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 2161.600 0.000 2162.160 0.560 ;
    END
  END caravel_io_pullup_sel[9]
  PIN caravel_io_schmitt_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 0.560 ;
    END
  END caravel_io_schmitt_sel[0]
  PIN caravel_io_schmitt_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2403.520 0.000 2404.080 0.560 ;
    END
  END caravel_io_schmitt_sel[10]
  PIN caravel_io_schmitt_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2618.560 0.000 2619.120 0.560 ;
    END
  END caravel_io_schmitt_sel[11]
  PIN caravel_io_schmitt_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2833.600 0.000 2834.160 0.560 ;
    END
  END caravel_io_schmitt_sel[12]
  PIN caravel_io_schmitt_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 0.560 ;
    END
  END caravel_io_schmitt_sel[1]
  PIN caravel_io_schmitt_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 0.560 ;
    END
  END caravel_io_schmitt_sel[2]
  PIN caravel_io_schmitt_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 898.240 0.000 898.800 0.560 ;
    END
  END caravel_io_schmitt_sel[3]
  PIN caravel_io_schmitt_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1113.280 0.000 1113.840 0.560 ;
    END
  END caravel_io_schmitt_sel[4]
  PIN caravel_io_schmitt_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1328.320 0.000 1328.880 0.560 ;
    END
  END caravel_io_schmitt_sel[5]
  PIN caravel_io_schmitt_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1543.360 0.000 1543.920 0.560 ;
    END
  END caravel_io_schmitt_sel[6]
  PIN caravel_io_schmitt_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1758.400 0.000 1758.960 0.560 ;
    END
  END caravel_io_schmitt_sel[7]
  PIN caravel_io_schmitt_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1973.440 0.000 1974.000 0.560 ;
    END
  END caravel_io_schmitt_sel[8]
  PIN caravel_io_schmitt_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2188.480 0.000 2189.040 0.560 ;
    END
  END caravel_io_schmitt_sel[9]
  PIN caravel_io_slew_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 0.560 ;
    END
  END caravel_io_slew_sel[0]
  PIN caravel_io_slew_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2430.400 0.000 2430.960 0.560 ;
    END
  END caravel_io_slew_sel[10]
  PIN caravel_io_slew_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2645.440 0.000 2646.000 0.560 ;
    END
  END caravel_io_slew_sel[11]
  PIN caravel_io_slew_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2860.480 0.000 2861.040 0.560 ;
    END
  END caravel_io_slew_sel[12]
  PIN caravel_io_slew_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 0.560 ;
    END
  END caravel_io_slew_sel[1]
  PIN caravel_io_slew_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 0.560 ;
    END
  END caravel_io_slew_sel[2]
  PIN caravel_io_slew_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 0.000 925.680 0.560 ;
    END
  END caravel_io_slew_sel[3]
  PIN caravel_io_slew_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1140.160 0.000 1140.720 0.560 ;
    END
  END caravel_io_slew_sel[4]
  PIN caravel_io_slew_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1355.200 0.000 1355.760 0.560 ;
    END
  END caravel_io_slew_sel[5]
  PIN caravel_io_slew_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1570.240 0.000 1570.800 0.560 ;
    END
  END caravel_io_slew_sel[6]
  PIN caravel_io_slew_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 1785.280 0.000 1785.840 0.560 ;
    END
  END caravel_io_slew_sel[7]
  PIN caravel_io_slew_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2000.320 0.000 2000.880 0.560 ;
    END
  END caravel_io_slew_sel[8]
  PIN caravel_io_slew_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2215.360 0.000 2215.920 0.560 ;
    END
  END caravel_io_slew_sel[9]
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.107000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 0.560 ;
    END
  END clock_core
  PIN flash_clk_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.130000 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 406.560 2900.000 407.120 ;
    END
  END flash_clk_frame
  PIN flash_clk_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 468.160 2900.000 468.720 ;
    END
  END flash_clk_oe
  PIN flash_csb_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.828000 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 283.360 2900.000 283.920 ;
    END
  END flash_csb_frame
  PIN flash_csb_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 344.960 2900.000 345.520 ;
    END
  END flash_csb_oe
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 529.760 2900.000 530.320 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.068800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 591.360 2900.000 591.920 ;
    END
  END flash_io0_do
  PIN flash_io0_ie
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.068800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 652.960 2900.000 653.520 ;
    END
  END flash_io0_ie
  PIN flash_io0_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.068800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 714.560 2900.000 715.120 ;
    END
  END flash_io0_oe
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 776.160 2900.000 776.720 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 837.760 2900.000 838.320 ;
    END
  END flash_io1_do
  PIN flash_io1_ie
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 899.360 2900.000 899.920 ;
    END
  END flash_io1_ie
  PIN flash_io1_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 960.960 2900.000 961.520 ;
    END
  END flash_io1_oe
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 36.960 2900.000 37.520 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 98.560 2900.000 99.120 ;
    END
  END gpio_inenb_core
  PIN gpio_out_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 160.160 2900.000 160.720 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal3 ;
        RECT 2899.440 221.760 2900.000 222.320 ;
    END
  END gpio_outenb_core
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 0.560 ;
    END
  END rstb
  PIN user_clock2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2096.640 999.440 2097.200 1000.000 ;
    END
  END user_clock2
  PIN user_gpio_in[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2115.680 999.440 2116.240 1000.000 ;
    END
  END user_gpio_in[0]
  PIN user_gpio_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2686.880 999.440 2687.440 1000.000 ;
    END
  END user_gpio_in[10]
  PIN user_gpio_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2744.000 999.440 2744.560 1000.000 ;
    END
  END user_gpio_in[11]
  PIN user_gpio_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2801.120 999.440 2801.680 1000.000 ;
    END
  END user_gpio_in[12]
  PIN user_gpio_in[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2172.800 999.440 2173.360 1000.000 ;
    END
  END user_gpio_in[1]
  PIN user_gpio_in[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal2 ;
        RECT 2229.920 999.440 2230.480 1000.000 ;
    END
  END user_gpio_in[2]
  PIN user_gpio_in[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2287.040 999.440 2287.600 1000.000 ;
    END
  END user_gpio_in[3]
  PIN user_gpio_in[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2344.160 999.440 2344.720 1000.000 ;
    END
  END user_gpio_in[4]
  PIN user_gpio_in[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2401.280 999.440 2401.840 1000.000 ;
    END
  END user_gpio_in[5]
  PIN user_gpio_in[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2458.400 999.440 2458.960 1000.000 ;
    END
  END user_gpio_in[6]
  PIN user_gpio_in[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2515.520 999.440 2516.080 1000.000 ;
    END
  END user_gpio_in[7]
  PIN user_gpio_in[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2572.640 999.440 2573.200 1000.000 ;
    END
  END user_gpio_in[8]
  PIN user_gpio_in[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2629.760 999.440 2630.320 1000.000 ;
    END
  END user_gpio_in[9]
  PIN user_gpio_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2134.720 999.440 2135.280 1000.000 ;
    END
  END user_gpio_oeb[0]
  PIN user_gpio_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2705.920 999.440 2706.480 1000.000 ;
    END
  END user_gpio_oeb[10]
  PIN user_gpio_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2763.040 999.440 2763.600 1000.000 ;
    END
  END user_gpio_oeb[11]
  PIN user_gpio_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2820.160 999.440 2820.720 1000.000 ;
    END
  END user_gpio_oeb[12]
  PIN user_gpio_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2191.840 999.440 2192.400 1000.000 ;
    END
  END user_gpio_oeb[1]
  PIN user_gpio_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 2248.960 999.440 2249.520 1000.000 ;
    END
  END user_gpio_oeb[2]
  PIN user_gpio_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 2306.080 999.440 2306.640 1000.000 ;
    END
  END user_gpio_oeb[3]
  PIN user_gpio_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2363.200 999.440 2363.760 1000.000 ;
    END
  END user_gpio_oeb[4]
  PIN user_gpio_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2420.320 999.440 2420.880 1000.000 ;
    END
  END user_gpio_oeb[5]
  PIN user_gpio_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2477.440 999.440 2478.000 1000.000 ;
    END
  END user_gpio_oeb[6]
  PIN user_gpio_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2534.560 999.440 2535.120 1000.000 ;
    END
  END user_gpio_oeb[7]
  PIN user_gpio_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2591.680 999.440 2592.240 1000.000 ;
    END
  END user_gpio_oeb[8]
  PIN user_gpio_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2648.800 999.440 2649.360 1000.000 ;
    END
  END user_gpio_oeb[9]
  PIN user_gpio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2153.760 999.440 2154.320 1000.000 ;
    END
  END user_gpio_out[0]
  PIN user_gpio_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2724.960 999.440 2725.520 1000.000 ;
    END
  END user_gpio_out[10]
  PIN user_gpio_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2782.080 999.440 2782.640 1000.000 ;
    END
  END user_gpio_out[11]
  PIN user_gpio_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2839.200 999.440 2839.760 1000.000 ;
    END
  END user_gpio_out[12]
  PIN user_gpio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2210.880 999.440 2211.440 1000.000 ;
    END
  END user_gpio_out[1]
  PIN user_gpio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 2268.000 999.440 2268.560 1000.000 ;
    END
  END user_gpio_out[2]
  PIN user_gpio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal2 ;
        RECT 2325.120 999.440 2325.680 1000.000 ;
    END
  END user_gpio_out[3]
  PIN user_gpio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2382.240 999.440 2382.800 1000.000 ;
    END
  END user_gpio_out[4]
  PIN user_gpio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2439.360 999.440 2439.920 1000.000 ;
    END
  END user_gpio_out[5]
  PIN user_gpio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2496.480 999.440 2497.040 1000.000 ;
    END
  END user_gpio_out[6]
  PIN user_gpio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2553.600 999.440 2554.160 1000.000 ;
    END
  END user_gpio_out[7]
  PIN user_gpio_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2610.720 999.440 2611.280 1000.000 ;
    END
  END user_gpio_out[8]
  PIN user_gpio_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 2667.840 999.440 2668.400 1000.000 ;
    END
  END user_gpio_out[9]
  PIN user_irq_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 2077.600 999.440 2078.160 1000.000 ;
    END
  END user_irq_core
  PIN user_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 999.440 2040.080 1000.000 ;
    END
  END user_wb_ack_i
  PIN user_wb_adr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 999.440 136.080 1000.000 ;
    END
  END user_wb_adr_o[0]
  PIN user_wb_adr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 999.440 326.480 1000.000 ;
    END
  END user_wb_adr_o[10]
  PIN user_wb_adr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 999.440 345.520 1000.000 ;
    END
  END user_wb_adr_o[11]
  PIN user_wb_adr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 999.440 364.560 1000.000 ;
    END
  END user_wb_adr_o[12]
  PIN user_wb_adr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 999.440 383.600 1000.000 ;
    END
  END user_wb_adr_o[13]
  PIN user_wb_adr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 999.440 402.640 1000.000 ;
    END
  END user_wb_adr_o[14]
  PIN user_wb_adr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 999.440 421.680 1000.000 ;
    END
  END user_wb_adr_o[15]
  PIN user_wb_adr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 999.440 440.720 1000.000 ;
    END
  END user_wb_adr_o[16]
  PIN user_wb_adr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 999.440 459.760 1000.000 ;
    END
  END user_wb_adr_o[17]
  PIN user_wb_adr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 999.440 478.800 1000.000 ;
    END
  END user_wb_adr_o[18]
  PIN user_wb_adr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 999.440 497.840 1000.000 ;
    END
  END user_wb_adr_o[19]
  PIN user_wb_adr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 999.440 155.120 1000.000 ;
    END
  END user_wb_adr_o[1]
  PIN user_wb_adr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 999.440 516.880 1000.000 ;
    END
  END user_wb_adr_o[20]
  PIN user_wb_adr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 999.440 535.920 1000.000 ;
    END
  END user_wb_adr_o[21]
  PIN user_wb_adr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 999.440 554.960 1000.000 ;
    END
  END user_wb_adr_o[22]
  PIN user_wb_adr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 573.440 999.440 574.000 1000.000 ;
    END
  END user_wb_adr_o[23]
  PIN user_wb_adr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 999.440 593.040 1000.000 ;
    END
  END user_wb_adr_o[24]
  PIN user_wb_adr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 999.440 612.080 1000.000 ;
    END
  END user_wb_adr_o[25]
  PIN user_wb_adr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 999.440 631.120 1000.000 ;
    END
  END user_wb_adr_o[26]
  PIN user_wb_adr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 999.440 650.160 1000.000 ;
    END
  END user_wb_adr_o[27]
  PIN user_wb_adr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 999.440 669.200 1000.000 ;
    END
  END user_wb_adr_o[28]
  PIN user_wb_adr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 999.440 688.240 1000.000 ;
    END
  END user_wb_adr_o[29]
  PIN user_wb_adr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 999.440 174.160 1000.000 ;
    END
  END user_wb_adr_o[2]
  PIN user_wb_adr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 999.440 707.280 1000.000 ;
    END
  END user_wb_adr_o[30]
  PIN user_wb_adr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 999.440 726.320 1000.000 ;
    END
  END user_wb_adr_o[31]
  PIN user_wb_adr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 999.440 193.200 1000.000 ;
    END
  END user_wb_adr_o[3]
  PIN user_wb_adr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 999.440 212.240 1000.000 ;
    END
  END user_wb_adr_o[4]
  PIN user_wb_adr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 999.440 231.280 1000.000 ;
    END
  END user_wb_adr_o[5]
  PIN user_wb_adr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 999.440 250.320 1000.000 ;
    END
  END user_wb_adr_o[6]
  PIN user_wb_adr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 999.440 269.360 1000.000 ;
    END
  END user_wb_adr_o[7]
  PIN user_wb_adr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 999.440 288.400 1000.000 ;
    END
  END user_wb_adr_o[8]
  PIN user_wb_adr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 999.440 307.440 1000.000 ;
    END
  END user_wb_adr_o[9]
  PIN user_wb_clk_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.130000 ;
    PORT
      LAYER Metal2 ;
        RECT 2058.560 999.440 2059.120 1000.000 ;
    END
  END user_wb_clk_o
  PIN user_wb_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1982.400 999.440 1982.960 1000.000 ;
    END
  END user_wb_cyc_o
  PIN user_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 999.440 1354.640 1000.000 ;
    END
  END user_wb_dat_i[0]
  PIN user_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1544.480 999.440 1545.040 1000.000 ;
    END
  END user_wb_dat_i[10]
  PIN user_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1563.520 999.440 1564.080 1000.000 ;
    END
  END user_wb_dat_i[11]
  PIN user_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 999.440 1583.120 1000.000 ;
    END
  END user_wb_dat_i[12]
  PIN user_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1601.600 999.440 1602.160 1000.000 ;
    END
  END user_wb_dat_i[13]
  PIN user_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1620.640 999.440 1621.200 1000.000 ;
    END
  END user_wb_dat_i[14]
  PIN user_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1639.680 999.440 1640.240 1000.000 ;
    END
  END user_wb_dat_i[15]
  PIN user_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1658.720 999.440 1659.280 1000.000 ;
    END
  END user_wb_dat_i[16]
  PIN user_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1677.760 999.440 1678.320 1000.000 ;
    END
  END user_wb_dat_i[17]
  PIN user_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 999.440 1697.360 1000.000 ;
    END
  END user_wb_dat_i[18]
  PIN user_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1715.840 999.440 1716.400 1000.000 ;
    END
  END user_wb_dat_i[19]
  PIN user_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1373.120 999.440 1373.680 1000.000 ;
    END
  END user_wb_dat_i[1]
  PIN user_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1734.880 999.440 1735.440 1000.000 ;
    END
  END user_wb_dat_i[20]
  PIN user_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1753.920 999.440 1754.480 1000.000 ;
    END
  END user_wb_dat_i[21]
  PIN user_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1772.960 999.440 1773.520 1000.000 ;
    END
  END user_wb_dat_i[22]
  PIN user_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1792.000 999.440 1792.560 1000.000 ;
    END
  END user_wb_dat_i[23]
  PIN user_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1811.040 999.440 1811.600 1000.000 ;
    END
  END user_wb_dat_i[24]
  PIN user_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1830.080 999.440 1830.640 1000.000 ;
    END
  END user_wb_dat_i[25]
  PIN user_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1849.120 999.440 1849.680 1000.000 ;
    END
  END user_wb_dat_i[26]
  PIN user_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1868.160 999.440 1868.720 1000.000 ;
    END
  END user_wb_dat_i[27]
  PIN user_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1887.200 999.440 1887.760 1000.000 ;
    END
  END user_wb_dat_i[28]
  PIN user_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 1906.240 999.440 1906.800 1000.000 ;
    END
  END user_wb_dat_i[29]
  PIN user_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 1392.160 999.440 1392.720 1000.000 ;
    END
  END user_wb_dat_i[2]
  PIN user_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 999.440 1925.840 1000.000 ;
    END
  END user_wb_dat_i[30]
  PIN user_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1944.320 999.440 1944.880 1000.000 ;
    END
  END user_wb_dat_i[31]
  PIN user_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 1411.200 999.440 1411.760 1000.000 ;
    END
  END user_wb_dat_i[3]
  PIN user_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1430.240 999.440 1430.800 1000.000 ;
    END
  END user_wb_dat_i[4]
  PIN user_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 1449.280 999.440 1449.840 1000.000 ;
    END
  END user_wb_dat_i[5]
  PIN user_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1468.320 999.440 1468.880 1000.000 ;
    END
  END user_wb_dat_i[6]
  PIN user_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1487.360 999.440 1487.920 1000.000 ;
    END
  END user_wb_dat_i[7]
  PIN user_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1506.400 999.440 1506.960 1000.000 ;
    END
  END user_wb_dat_i[8]
  PIN user_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal2 ;
        RECT 1525.440 999.440 1526.000 1000.000 ;
    END
  END user_wb_dat_i[9]
  PIN user_wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 744.800 999.440 745.360 1000.000 ;
    END
  END user_wb_dat_o[0]
  PIN user_wb_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 999.440 935.760 1000.000 ;
    END
  END user_wb_dat_o[10]
  PIN user_wb_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 999.440 954.800 1000.000 ;
    END
  END user_wb_dat_o[11]
  PIN user_wb_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 999.440 973.840 1000.000 ;
    END
  END user_wb_dat_o[12]
  PIN user_wb_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 992.320 999.440 992.880 1000.000 ;
    END
  END user_wb_dat_o[13]
  PIN user_wb_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 999.440 1011.920 1000.000 ;
    END
  END user_wb_dat_o[14]
  PIN user_wb_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1030.400 999.440 1030.960 1000.000 ;
    END
  END user_wb_dat_o[15]
  PIN user_wb_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1049.440 999.440 1050.000 1000.000 ;
    END
  END user_wb_dat_o[16]
  PIN user_wb_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 999.440 1069.040 1000.000 ;
    END
  END user_wb_dat_o[17]
  PIN user_wb_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1087.520 999.440 1088.080 1000.000 ;
    END
  END user_wb_dat_o[18]
  PIN user_wb_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1106.560 999.440 1107.120 1000.000 ;
    END
  END user_wb_dat_o[19]
  PIN user_wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 999.440 764.400 1000.000 ;
    END
  END user_wb_dat_o[1]
  PIN user_wb_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 999.440 1126.160 1000.000 ;
    END
  END user_wb_dat_o[20]
  PIN user_wb_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1144.640 999.440 1145.200 1000.000 ;
    END
  END user_wb_dat_o[21]
  PIN user_wb_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1163.680 999.440 1164.240 1000.000 ;
    END
  END user_wb_dat_o[22]
  PIN user_wb_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1182.720 999.440 1183.280 1000.000 ;
    END
  END user_wb_dat_o[23]
  PIN user_wb_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1201.760 999.440 1202.320 1000.000 ;
    END
  END user_wb_dat_o[24]
  PIN user_wb_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1220.800 999.440 1221.360 1000.000 ;
    END
  END user_wb_dat_o[25]
  PIN user_wb_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1239.840 999.440 1240.400 1000.000 ;
    END
  END user_wb_dat_o[26]
  PIN user_wb_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1258.880 999.440 1259.440 1000.000 ;
    END
  END user_wb_dat_o[27]
  PIN user_wb_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1277.920 999.440 1278.480 1000.000 ;
    END
  END user_wb_dat_o[28]
  PIN user_wb_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1296.960 999.440 1297.520 1000.000 ;
    END
  END user_wb_dat_o[29]
  PIN user_wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 999.440 783.440 1000.000 ;
    END
  END user_wb_dat_o[2]
  PIN user_wb_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1316.000 999.440 1316.560 1000.000 ;
    END
  END user_wb_dat_o[30]
  PIN user_wb_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1335.040 999.440 1335.600 1000.000 ;
    END
  END user_wb_dat_o[31]
  PIN user_wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 999.440 802.480 1000.000 ;
    END
  END user_wb_dat_o[3]
  PIN user_wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 999.440 821.520 1000.000 ;
    END
  END user_wb_dat_o[4]
  PIN user_wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 999.440 840.560 1000.000 ;
    END
  END user_wb_dat_o[5]
  PIN user_wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 859.040 999.440 859.600 1000.000 ;
    END
  END user_wb_dat_o[6]
  PIN user_wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 999.440 878.640 1000.000 ;
    END
  END user_wb_dat_o[7]
  PIN user_wb_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 999.440 897.680 1000.000 ;
    END
  END user_wb_dat_o[8]
  PIN user_wb_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 999.440 916.720 1000.000 ;
    END
  END user_wb_dat_o[9]
  PIN user_wb_rst_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 1963.360 999.440 1963.920 1000.000 ;
    END
  END user_wb_rst_o
  PIN user_wb_sel_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 999.440 59.920 1000.000 ;
    END
  END user_wb_sel_o[0]
  PIN user_wb_sel_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 999.440 78.960 1000.000 ;
    END
  END user_wb_sel_o[1]
  PIN user_wb_sel_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 999.440 98.000 1000.000 ;
    END
  END user_wb_sel_o[2]
  PIN user_wb_sel_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 999.440 117.040 1000.000 ;
    END
  END user_wb_sel_o[3]
  PIN user_wb_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2001.440 999.440 2002.000 1000.000 ;
    END
  END user_wb_stb_o
  PIN user_wb_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal2 ;
        RECT 2020.480 999.440 2021.040 1000.000 ;
    END
  END user_wb_we_o
  OBS
      LAYER Nwell ;
        RECT 23.650 27.010 2874.910 972.590 ;
      LAYER Metal1 ;
        RECT 24.080 27.140 2874.480 972.460 ;
      LAYER Metal2 ;
        RECT 25.340 999.140 59.060 999.860 ;
        RECT 60.220 999.140 78.100 999.860 ;
        RECT 79.260 999.140 97.140 999.860 ;
        RECT 98.300 999.140 116.180 999.860 ;
        RECT 117.340 999.140 135.220 999.860 ;
        RECT 136.380 999.140 154.260 999.860 ;
        RECT 155.420 999.140 173.300 999.860 ;
        RECT 174.460 999.140 192.340 999.860 ;
        RECT 193.500 999.140 211.380 999.860 ;
        RECT 212.540 999.140 230.420 999.860 ;
        RECT 231.580 999.140 249.460 999.860 ;
        RECT 250.620 999.140 268.500 999.860 ;
        RECT 269.660 999.140 287.540 999.860 ;
        RECT 288.700 999.140 306.580 999.860 ;
        RECT 307.740 999.140 325.620 999.860 ;
        RECT 326.780 999.140 344.660 999.860 ;
        RECT 345.820 999.140 363.700 999.860 ;
        RECT 364.860 999.140 382.740 999.860 ;
        RECT 383.900 999.140 401.780 999.860 ;
        RECT 402.940 999.140 420.820 999.860 ;
        RECT 421.980 999.140 439.860 999.860 ;
        RECT 441.020 999.140 458.900 999.860 ;
        RECT 460.060 999.140 477.940 999.860 ;
        RECT 479.100 999.140 496.980 999.860 ;
        RECT 498.140 999.140 516.020 999.860 ;
        RECT 517.180 999.140 535.060 999.860 ;
        RECT 536.220 999.140 554.100 999.860 ;
        RECT 555.260 999.140 573.140 999.860 ;
        RECT 574.300 999.140 592.180 999.860 ;
        RECT 593.340 999.140 611.220 999.860 ;
        RECT 612.380 999.140 630.260 999.860 ;
        RECT 631.420 999.140 649.300 999.860 ;
        RECT 650.460 999.140 668.340 999.860 ;
        RECT 669.500 999.140 687.380 999.860 ;
        RECT 688.540 999.140 706.420 999.860 ;
        RECT 707.580 999.140 725.460 999.860 ;
        RECT 726.620 999.140 744.500 999.860 ;
        RECT 745.660 999.140 763.540 999.860 ;
        RECT 764.700 999.140 782.580 999.860 ;
        RECT 783.740 999.140 801.620 999.860 ;
        RECT 802.780 999.140 820.660 999.860 ;
        RECT 821.820 999.140 839.700 999.860 ;
        RECT 840.860 999.140 858.740 999.860 ;
        RECT 859.900 999.140 877.780 999.860 ;
        RECT 878.940 999.140 896.820 999.860 ;
        RECT 897.980 999.140 915.860 999.860 ;
        RECT 917.020 999.140 934.900 999.860 ;
        RECT 936.060 999.140 953.940 999.860 ;
        RECT 955.100 999.140 972.980 999.860 ;
        RECT 974.140 999.140 992.020 999.860 ;
        RECT 993.180 999.140 1011.060 999.860 ;
        RECT 1012.220 999.140 1030.100 999.860 ;
        RECT 1031.260 999.140 1049.140 999.860 ;
        RECT 1050.300 999.140 1068.180 999.860 ;
        RECT 1069.340 999.140 1087.220 999.860 ;
        RECT 1088.380 999.140 1106.260 999.860 ;
        RECT 1107.420 999.140 1125.300 999.860 ;
        RECT 1126.460 999.140 1144.340 999.860 ;
        RECT 1145.500 999.140 1163.380 999.860 ;
        RECT 1164.540 999.140 1182.420 999.860 ;
        RECT 1183.580 999.140 1201.460 999.860 ;
        RECT 1202.620 999.140 1220.500 999.860 ;
        RECT 1221.660 999.140 1239.540 999.860 ;
        RECT 1240.700 999.140 1258.580 999.860 ;
        RECT 1259.740 999.140 1277.620 999.860 ;
        RECT 1278.780 999.140 1296.660 999.860 ;
        RECT 1297.820 999.140 1315.700 999.860 ;
        RECT 1316.860 999.140 1334.740 999.860 ;
        RECT 1335.900 999.140 1353.780 999.860 ;
        RECT 1354.940 999.140 1372.820 999.860 ;
        RECT 1373.980 999.140 1391.860 999.860 ;
        RECT 1393.020 999.140 1410.900 999.860 ;
        RECT 1412.060 999.140 1429.940 999.860 ;
        RECT 1431.100 999.140 1448.980 999.860 ;
        RECT 1450.140 999.140 1468.020 999.860 ;
        RECT 1469.180 999.140 1487.060 999.860 ;
        RECT 1488.220 999.140 1506.100 999.860 ;
        RECT 1507.260 999.140 1525.140 999.860 ;
        RECT 1526.300 999.140 1544.180 999.860 ;
        RECT 1545.340 999.140 1563.220 999.860 ;
        RECT 1564.380 999.140 1582.260 999.860 ;
        RECT 1583.420 999.140 1601.300 999.860 ;
        RECT 1602.460 999.140 1620.340 999.860 ;
        RECT 1621.500 999.140 1639.380 999.860 ;
        RECT 1640.540 999.140 1658.420 999.860 ;
        RECT 1659.580 999.140 1677.460 999.860 ;
        RECT 1678.620 999.140 1696.500 999.860 ;
        RECT 1697.660 999.140 1715.540 999.860 ;
        RECT 1716.700 999.140 1734.580 999.860 ;
        RECT 1735.740 999.140 1753.620 999.860 ;
        RECT 1754.780 999.140 1772.660 999.860 ;
        RECT 1773.820 999.140 1791.700 999.860 ;
        RECT 1792.860 999.140 1810.740 999.860 ;
        RECT 1811.900 999.140 1829.780 999.860 ;
        RECT 1830.940 999.140 1848.820 999.860 ;
        RECT 1849.980 999.140 1867.860 999.860 ;
        RECT 1869.020 999.140 1886.900 999.860 ;
        RECT 1888.060 999.140 1905.940 999.860 ;
        RECT 1907.100 999.140 1924.980 999.860 ;
        RECT 1926.140 999.140 1944.020 999.860 ;
        RECT 1945.180 999.140 1963.060 999.860 ;
        RECT 1964.220 999.140 1982.100 999.860 ;
        RECT 1983.260 999.140 2001.140 999.860 ;
        RECT 2002.300 999.140 2020.180 999.860 ;
        RECT 2021.340 999.140 2039.220 999.860 ;
        RECT 2040.380 999.140 2058.260 999.860 ;
        RECT 2059.420 999.140 2077.300 999.860 ;
        RECT 2078.460 999.140 2096.340 999.860 ;
        RECT 2097.500 999.140 2115.380 999.860 ;
        RECT 2116.540 999.140 2134.420 999.860 ;
        RECT 2135.580 999.140 2153.460 999.860 ;
        RECT 2154.620 999.140 2172.500 999.860 ;
        RECT 2173.660 999.140 2191.540 999.860 ;
        RECT 2192.700 999.140 2210.580 999.860 ;
        RECT 2211.740 999.140 2229.620 999.860 ;
        RECT 2230.780 999.140 2248.660 999.860 ;
        RECT 2249.820 999.140 2267.700 999.860 ;
        RECT 2268.860 999.140 2286.740 999.860 ;
        RECT 2287.900 999.140 2305.780 999.860 ;
        RECT 2306.940 999.140 2324.820 999.860 ;
        RECT 2325.980 999.140 2343.860 999.860 ;
        RECT 2345.020 999.140 2362.900 999.860 ;
        RECT 2364.060 999.140 2381.940 999.860 ;
        RECT 2383.100 999.140 2400.980 999.860 ;
        RECT 2402.140 999.140 2420.020 999.860 ;
        RECT 2421.180 999.140 2439.060 999.860 ;
        RECT 2440.220 999.140 2458.100 999.860 ;
        RECT 2459.260 999.140 2477.140 999.860 ;
        RECT 2478.300 999.140 2496.180 999.860 ;
        RECT 2497.340 999.140 2515.220 999.860 ;
        RECT 2516.380 999.140 2534.260 999.860 ;
        RECT 2535.420 999.140 2553.300 999.860 ;
        RECT 2554.460 999.140 2572.340 999.860 ;
        RECT 2573.500 999.140 2591.380 999.860 ;
        RECT 2592.540 999.140 2610.420 999.860 ;
        RECT 2611.580 999.140 2629.460 999.860 ;
        RECT 2630.620 999.140 2648.500 999.860 ;
        RECT 2649.660 999.140 2667.540 999.860 ;
        RECT 2668.700 999.140 2686.580 999.860 ;
        RECT 2687.740 999.140 2705.620 999.860 ;
        RECT 2706.780 999.140 2724.660 999.860 ;
        RECT 2725.820 999.140 2743.700 999.860 ;
        RECT 2744.860 999.140 2762.740 999.860 ;
        RECT 2763.900 999.140 2781.780 999.860 ;
        RECT 2782.940 999.140 2800.820 999.860 ;
        RECT 2801.980 999.140 2819.860 999.860 ;
        RECT 2821.020 999.140 2838.900 999.860 ;
        RECT 2840.060 999.140 2872.660 999.860 ;
        RECT 25.340 0.860 2872.660 999.140 ;
        RECT 25.340 0.090 37.780 0.860 ;
        RECT 38.940 0.090 64.660 0.860 ;
        RECT 65.820 0.090 91.540 0.860 ;
        RECT 92.700 0.090 118.420 0.860 ;
        RECT 119.580 0.090 145.300 0.860 ;
        RECT 146.460 0.090 172.180 0.860 ;
        RECT 173.340 0.090 199.060 0.860 ;
        RECT 200.220 0.090 225.940 0.860 ;
        RECT 227.100 0.090 252.820 0.860 ;
        RECT 253.980 0.090 279.700 0.860 ;
        RECT 280.860 0.090 306.580 0.860 ;
        RECT 307.740 0.090 333.460 0.860 ;
        RECT 334.620 0.090 360.340 0.860 ;
        RECT 361.500 0.090 387.220 0.860 ;
        RECT 388.380 0.090 414.100 0.860 ;
        RECT 415.260 0.090 440.980 0.860 ;
        RECT 442.140 0.090 467.860 0.860 ;
        RECT 469.020 0.090 494.740 0.860 ;
        RECT 495.900 0.090 521.620 0.860 ;
        RECT 522.780 0.090 548.500 0.860 ;
        RECT 549.660 0.090 575.380 0.860 ;
        RECT 576.540 0.090 602.260 0.860 ;
        RECT 603.420 0.090 629.140 0.860 ;
        RECT 630.300 0.090 656.020 0.860 ;
        RECT 657.180 0.090 682.900 0.860 ;
        RECT 684.060 0.090 709.780 0.860 ;
        RECT 710.940 0.090 736.660 0.860 ;
        RECT 737.820 0.090 763.540 0.860 ;
        RECT 764.700 0.090 790.420 0.860 ;
        RECT 791.580 0.090 817.300 0.860 ;
        RECT 818.460 0.090 844.180 0.860 ;
        RECT 845.340 0.090 871.060 0.860 ;
        RECT 872.220 0.090 897.940 0.860 ;
        RECT 899.100 0.090 924.820 0.860 ;
        RECT 925.980 0.090 951.700 0.860 ;
        RECT 952.860 0.090 978.580 0.860 ;
        RECT 979.740 0.090 1005.460 0.860 ;
        RECT 1006.620 0.090 1032.340 0.860 ;
        RECT 1033.500 0.090 1059.220 0.860 ;
        RECT 1060.380 0.090 1086.100 0.860 ;
        RECT 1087.260 0.090 1112.980 0.860 ;
        RECT 1114.140 0.090 1139.860 0.860 ;
        RECT 1141.020 0.090 1166.740 0.860 ;
        RECT 1167.900 0.090 1193.620 0.860 ;
        RECT 1194.780 0.090 1220.500 0.860 ;
        RECT 1221.660 0.090 1247.380 0.860 ;
        RECT 1248.540 0.090 1274.260 0.860 ;
        RECT 1275.420 0.090 1301.140 0.860 ;
        RECT 1302.300 0.090 1328.020 0.860 ;
        RECT 1329.180 0.090 1354.900 0.860 ;
        RECT 1356.060 0.090 1381.780 0.860 ;
        RECT 1382.940 0.090 1408.660 0.860 ;
        RECT 1409.820 0.090 1435.540 0.860 ;
        RECT 1436.700 0.090 1462.420 0.860 ;
        RECT 1463.580 0.090 1489.300 0.860 ;
        RECT 1490.460 0.090 1516.180 0.860 ;
        RECT 1517.340 0.090 1543.060 0.860 ;
        RECT 1544.220 0.090 1569.940 0.860 ;
        RECT 1571.100 0.090 1596.820 0.860 ;
        RECT 1597.980 0.090 1623.700 0.860 ;
        RECT 1624.860 0.090 1650.580 0.860 ;
        RECT 1651.740 0.090 1677.460 0.860 ;
        RECT 1678.620 0.090 1704.340 0.860 ;
        RECT 1705.500 0.090 1731.220 0.860 ;
        RECT 1732.380 0.090 1758.100 0.860 ;
        RECT 1759.260 0.090 1784.980 0.860 ;
        RECT 1786.140 0.090 1811.860 0.860 ;
        RECT 1813.020 0.090 1838.740 0.860 ;
        RECT 1839.900 0.090 1865.620 0.860 ;
        RECT 1866.780 0.090 1892.500 0.860 ;
        RECT 1893.660 0.090 1919.380 0.860 ;
        RECT 1920.540 0.090 1946.260 0.860 ;
        RECT 1947.420 0.090 1973.140 0.860 ;
        RECT 1974.300 0.090 2000.020 0.860 ;
        RECT 2001.180 0.090 2026.900 0.860 ;
        RECT 2028.060 0.090 2053.780 0.860 ;
        RECT 2054.940 0.090 2080.660 0.860 ;
        RECT 2081.820 0.090 2107.540 0.860 ;
        RECT 2108.700 0.090 2134.420 0.860 ;
        RECT 2135.580 0.090 2161.300 0.860 ;
        RECT 2162.460 0.090 2188.180 0.860 ;
        RECT 2189.340 0.090 2215.060 0.860 ;
        RECT 2216.220 0.090 2241.940 0.860 ;
        RECT 2243.100 0.090 2268.820 0.860 ;
        RECT 2269.980 0.090 2295.700 0.860 ;
        RECT 2296.860 0.090 2322.580 0.860 ;
        RECT 2323.740 0.090 2349.460 0.860 ;
        RECT 2350.620 0.090 2376.340 0.860 ;
        RECT 2377.500 0.090 2403.220 0.860 ;
        RECT 2404.380 0.090 2430.100 0.860 ;
        RECT 2431.260 0.090 2456.980 0.860 ;
        RECT 2458.140 0.090 2483.860 0.860 ;
        RECT 2485.020 0.090 2510.740 0.860 ;
        RECT 2511.900 0.090 2537.620 0.860 ;
        RECT 2538.780 0.090 2564.500 0.860 ;
        RECT 2565.660 0.090 2591.380 0.860 ;
        RECT 2592.540 0.090 2618.260 0.860 ;
        RECT 2619.420 0.090 2645.140 0.860 ;
        RECT 2646.300 0.090 2672.020 0.860 ;
        RECT 2673.180 0.090 2698.900 0.860 ;
        RECT 2700.060 0.090 2725.780 0.860 ;
        RECT 2726.940 0.090 2752.660 0.860 ;
        RECT 2753.820 0.090 2779.540 0.860 ;
        RECT 2780.700 0.090 2806.420 0.860 ;
        RECT 2807.580 0.090 2833.300 0.860 ;
        RECT 2834.460 0.090 2860.180 0.860 ;
        RECT 2861.340 0.090 2872.660 0.860 ;
      LAYER Metal3 ;
        RECT 25.290 961.820 2899.440 999.460 ;
        RECT 25.290 960.660 2899.140 961.820 ;
        RECT 25.290 900.220 2899.440 960.660 ;
        RECT 25.290 899.060 2899.140 900.220 ;
        RECT 25.290 838.620 2899.440 899.060 ;
        RECT 25.290 837.460 2899.140 838.620 ;
        RECT 25.290 777.020 2899.440 837.460 ;
        RECT 25.290 775.860 2899.140 777.020 ;
        RECT 25.290 715.420 2899.440 775.860 ;
        RECT 25.290 714.260 2899.140 715.420 ;
        RECT 25.290 653.820 2899.440 714.260 ;
        RECT 25.290 652.660 2899.140 653.820 ;
        RECT 25.290 592.220 2899.440 652.660 ;
        RECT 25.290 591.060 2899.140 592.220 ;
        RECT 25.290 530.620 2899.440 591.060 ;
        RECT 25.290 529.460 2899.140 530.620 ;
        RECT 25.290 469.020 2899.440 529.460 ;
        RECT 25.290 467.860 2899.140 469.020 ;
        RECT 25.290 407.420 2899.440 467.860 ;
        RECT 25.290 406.260 2899.140 407.420 ;
        RECT 25.290 345.820 2899.440 406.260 ;
        RECT 25.290 344.660 2899.140 345.820 ;
        RECT 25.290 284.220 2899.440 344.660 ;
        RECT 25.290 283.060 2899.140 284.220 ;
        RECT 25.290 222.620 2899.440 283.060 ;
        RECT 25.290 221.460 2899.140 222.620 ;
        RECT 25.290 161.020 2899.440 221.460 ;
        RECT 25.290 159.860 2899.140 161.020 ;
        RECT 25.290 99.420 2899.440 159.860 ;
        RECT 25.290 98.260 2899.140 99.420 ;
        RECT 25.290 37.820 2899.440 98.260 ;
        RECT 25.290 36.660 2899.140 37.820 ;
        RECT 25.290 0.140 2899.440 36.660 ;
      LAYER Metal4 ;
        RECT 46.620 994.460 2851.940 997.830 ;
        RECT 46.620 5.140 47.780 994.460 ;
        RECT 51.380 5.140 105.780 994.460 ;
        RECT 109.380 5.140 127.780 994.460 ;
        RECT 131.380 5.140 185.780 994.460 ;
        RECT 189.380 5.140 207.780 994.460 ;
        RECT 211.380 5.140 265.780 994.460 ;
        RECT 269.380 5.140 287.780 994.460 ;
        RECT 291.380 5.140 345.780 994.460 ;
        RECT 349.380 5.140 367.780 994.460 ;
        RECT 371.380 5.140 425.780 994.460 ;
        RECT 429.380 5.140 447.780 994.460 ;
        RECT 451.380 5.140 505.780 994.460 ;
        RECT 509.380 5.140 527.780 994.460 ;
        RECT 531.380 5.140 585.780 994.460 ;
        RECT 589.380 5.140 607.780 994.460 ;
        RECT 611.380 545.500 665.780 994.460 ;
        RECT 669.380 545.500 687.780 994.460 ;
        RECT 611.380 66.420 687.780 545.500 ;
        RECT 611.380 5.140 665.780 66.420 ;
        RECT 669.380 5.140 687.780 66.420 ;
        RECT 691.380 5.140 745.780 994.460 ;
        RECT 749.380 5.140 767.780 994.460 ;
        RECT 771.380 5.140 825.780 994.460 ;
        RECT 829.380 5.140 847.780 994.460 ;
        RECT 851.380 5.140 905.780 994.460 ;
        RECT 909.380 5.140 927.780 994.460 ;
        RECT 931.380 5.140 985.780 994.460 ;
        RECT 989.380 5.140 1007.780 994.460 ;
        RECT 1011.380 5.140 1065.780 994.460 ;
        RECT 1069.380 545.500 1087.780 994.460 ;
        RECT 1091.380 545.500 1145.780 994.460 ;
        RECT 1069.380 66.420 1145.780 545.500 ;
        RECT 1069.380 5.140 1087.780 66.420 ;
        RECT 1091.380 5.140 1145.780 66.420 ;
        RECT 1149.380 5.140 1167.780 994.460 ;
        RECT 1171.380 5.140 1225.780 994.460 ;
        RECT 1229.380 5.140 1247.780 994.460 ;
        RECT 1251.380 5.140 1305.780 994.460 ;
        RECT 1309.380 5.140 1327.780 994.460 ;
        RECT 1331.380 5.140 1385.780 994.460 ;
        RECT 1389.380 5.140 1407.780 994.460 ;
        RECT 1411.380 5.140 1465.780 994.460 ;
        RECT 1469.380 5.140 1487.780 994.460 ;
        RECT 1491.380 5.140 1545.780 994.460 ;
        RECT 1549.380 5.140 1567.780 994.460 ;
        RECT 1571.380 5.140 1625.780 994.460 ;
        RECT 1629.380 5.140 1647.780 994.460 ;
        RECT 1651.380 5.140 1705.780 994.460 ;
        RECT 1709.380 5.140 1727.780 994.460 ;
        RECT 1731.380 5.140 1785.780 994.460 ;
        RECT 1789.380 5.140 1807.780 994.460 ;
        RECT 1811.380 5.140 1865.780 994.460 ;
        RECT 1869.380 5.140 1887.780 994.460 ;
        RECT 1891.380 5.140 1945.780 994.460 ;
        RECT 1949.380 5.140 1967.780 994.460 ;
        RECT 1971.380 5.140 2025.780 994.460 ;
        RECT 2029.380 5.140 2047.780 994.460 ;
        RECT 2051.380 5.140 2105.780 994.460 ;
        RECT 2109.380 5.140 2127.780 994.460 ;
        RECT 2131.380 5.140 2185.780 994.460 ;
        RECT 2189.380 5.140 2207.780 994.460 ;
        RECT 2211.380 5.140 2265.780 994.460 ;
        RECT 2269.380 5.140 2287.780 994.460 ;
        RECT 2291.380 5.140 2345.780 994.460 ;
        RECT 2349.380 5.140 2367.780 994.460 ;
        RECT 2371.380 5.140 2425.780 994.460 ;
        RECT 2429.380 5.140 2447.780 994.460 ;
        RECT 2451.380 5.140 2505.780 994.460 ;
        RECT 2509.380 5.140 2527.780 994.460 ;
        RECT 2531.380 5.140 2585.780 994.460 ;
        RECT 2589.380 5.140 2607.780 994.460 ;
        RECT 2611.380 5.140 2620.280 994.460 ;
        RECT 2623.880 5.140 2632.280 994.460 ;
        RECT 2635.880 144.425 2665.780 994.460 ;
        RECT 2669.380 144.425 2687.780 994.460 ;
        RECT 2691.380 144.425 2745.780 994.460 ;
        RECT 2635.880 87.030 2745.780 144.425 ;
        RECT 2635.880 5.140 2665.780 87.030 ;
        RECT 2669.380 5.140 2687.780 87.030 ;
        RECT 2691.380 5.140 2745.780 87.030 ;
        RECT 2749.380 5.140 2767.780 994.460 ;
        RECT 2771.380 5.140 2825.780 994.460 ;
        RECT 2829.380 5.140 2847.780 994.460 ;
        RECT 2851.380 5.140 2851.940 994.460 ;
        RECT 46.620 1.210 2851.940 5.140 ;
      LAYER Metal5 ;
        RECT 63.340 994.760 2830.740 996.970 ;
        RECT 63.340 982.760 2830.740 983.560 ;
        RECT 63.340 960.190 2830.740 971.560 ;
        RECT 63.340 930.190 2830.740 955.990 ;
        RECT 63.340 900.190 2830.740 925.990 ;
        RECT 63.340 870.190 2830.740 895.990 ;
        RECT 63.340 840.190 2830.740 865.990 ;
        RECT 63.340 810.190 2830.740 835.990 ;
        RECT 63.340 780.190 2830.740 805.990 ;
        RECT 63.340 750.190 2830.740 775.990 ;
        RECT 63.340 720.190 2830.740 745.990 ;
        RECT 63.340 690.190 2830.740 715.990 ;
        RECT 63.340 660.190 2830.740 685.990 ;
        RECT 63.340 630.190 2830.740 655.990 ;
        RECT 63.340 600.190 2830.740 625.990 ;
        RECT 63.340 570.190 2830.740 595.990 ;
        RECT 63.340 540.190 2830.740 565.990 ;
        RECT 63.340 510.190 2830.740 535.990 ;
        RECT 63.340 480.190 2830.740 505.990 ;
        RECT 63.340 450.190 2830.740 475.990 ;
        RECT 63.340 420.190 2830.740 445.990 ;
        RECT 63.340 390.190 2830.740 415.990 ;
        RECT 63.340 360.190 2830.740 385.990 ;
        RECT 63.340 330.190 2830.740 355.990 ;
        RECT 63.340 300.190 2830.740 325.990 ;
        RECT 63.340 270.190 2830.740 295.990 ;
        RECT 63.340 240.190 2830.740 265.990 ;
        RECT 63.340 210.190 2830.740 235.990 ;
        RECT 63.340 180.190 2830.740 205.990 ;
        RECT 63.340 150.190 2830.740 175.990 ;
        RECT 2636.495 145.990 2706.855 150.190 ;
        RECT 63.340 120.190 2830.740 145.990 ;
        RECT 2636.495 115.990 2706.855 120.190 ;
        RECT 63.340 90.190 2830.740 115.990 ;
        RECT 2636.995 85.990 2706.855 90.190 ;
        RECT 63.340 60.190 2830.740 85.990 ;
        RECT 63.340 32.630 2830.740 55.990 ;
  END
END caravel_core
END LIBRARY

