module efuse_wb_mem_128x8 (wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rst_i,
    wb_sel_i,
    wb_stb_i,
    wb_we_i,
    write_enable_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o);
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rst_i;
 input wb_sel_i;
 input wb_stb_i;
 input wb_we_i;
 input write_enable_i;
 input [6:0] wb_adr_i;
 input [7:0] wb_dat_i;
 output [7:0] wb_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire \bit_sel[0] ;
 wire \bit_sel[10] ;
 wire \bit_sel[11] ;
 wire \bit_sel[12] ;
 wire \bit_sel[13] ;
 wire \bit_sel[14] ;
 wire \bit_sel[15] ;
 wire \bit_sel[16] ;
 wire \bit_sel[17] ;
 wire \bit_sel[18] ;
 wire \bit_sel[19] ;
 wire \bit_sel[1] ;
 wire \bit_sel[20] ;
 wire \bit_sel[21] ;
 wire \bit_sel[22] ;
 wire \bit_sel[23] ;
 wire \bit_sel[24] ;
 wire \bit_sel[25] ;
 wire \bit_sel[26] ;
 wire \bit_sel[27] ;
 wire \bit_sel[28] ;
 wire \bit_sel[29] ;
 wire \bit_sel[2] ;
 wire \bit_sel[30] ;
 wire \bit_sel[31] ;
 wire \bit_sel[32] ;
 wire \bit_sel[33] ;
 wire \bit_sel[34] ;
 wire \bit_sel[35] ;
 wire \bit_sel[36] ;
 wire \bit_sel[37] ;
 wire \bit_sel[38] ;
 wire \bit_sel[39] ;
 wire \bit_sel[3] ;
 wire \bit_sel[40] ;
 wire \bit_sel[41] ;
 wire \bit_sel[42] ;
 wire \bit_sel[43] ;
 wire \bit_sel[44] ;
 wire \bit_sel[45] ;
 wire \bit_sel[46] ;
 wire \bit_sel[47] ;
 wire \bit_sel[48] ;
 wire \bit_sel[49] ;
 wire \bit_sel[4] ;
 wire \bit_sel[50] ;
 wire \bit_sel[51] ;
 wire \bit_sel[52] ;
 wire \bit_sel[53] ;
 wire \bit_sel[54] ;
 wire \bit_sel[55] ;
 wire \bit_sel[56] ;
 wire \bit_sel[57] ;
 wire \bit_sel[58] ;
 wire \bit_sel[59] ;
 wire \bit_sel[5] ;
 wire \bit_sel[60] ;
 wire \bit_sel[61] ;
 wire \bit_sel[62] ;
 wire \bit_sel[63] ;
 wire \bit_sel[6] ;
 wire \bit_sel[7] ;
 wire \bit_sel[8] ;
 wire \bit_sel[9] ;
 wire \bit_sel_reg[0] ;
 wire \bit_sel_reg[10] ;
 wire \bit_sel_reg[11] ;
 wire \bit_sel_reg[12] ;
 wire \bit_sel_reg[13] ;
 wire \bit_sel_reg[14] ;
 wire \bit_sel_reg[15] ;
 wire \bit_sel_reg[16] ;
 wire \bit_sel_reg[17] ;
 wire \bit_sel_reg[18] ;
 wire \bit_sel_reg[19] ;
 wire \bit_sel_reg[1] ;
 wire \bit_sel_reg[20] ;
 wire \bit_sel_reg[21] ;
 wire \bit_sel_reg[22] ;
 wire \bit_sel_reg[23] ;
 wire \bit_sel_reg[24] ;
 wire \bit_sel_reg[25] ;
 wire \bit_sel_reg[26] ;
 wire \bit_sel_reg[27] ;
 wire \bit_sel_reg[28] ;
 wire \bit_sel_reg[29] ;
 wire \bit_sel_reg[2] ;
 wire \bit_sel_reg[30] ;
 wire \bit_sel_reg[31] ;
 wire \bit_sel_reg[32] ;
 wire \bit_sel_reg[33] ;
 wire \bit_sel_reg[34] ;
 wire \bit_sel_reg[35] ;
 wire \bit_sel_reg[36] ;
 wire \bit_sel_reg[37] ;
 wire \bit_sel_reg[38] ;
 wire \bit_sel_reg[39] ;
 wire \bit_sel_reg[3] ;
 wire \bit_sel_reg[40] ;
 wire \bit_sel_reg[41] ;
 wire \bit_sel_reg[42] ;
 wire \bit_sel_reg[43] ;
 wire \bit_sel_reg[44] ;
 wire \bit_sel_reg[45] ;
 wire \bit_sel_reg[46] ;
 wire \bit_sel_reg[47] ;
 wire \bit_sel_reg[48] ;
 wire \bit_sel_reg[49] ;
 wire \bit_sel_reg[4] ;
 wire \bit_sel_reg[50] ;
 wire \bit_sel_reg[51] ;
 wire \bit_sel_reg[52] ;
 wire \bit_sel_reg[53] ;
 wire \bit_sel_reg[54] ;
 wire \bit_sel_reg[55] ;
 wire \bit_sel_reg[56] ;
 wire \bit_sel_reg[57] ;
 wire \bit_sel_reg[58] ;
 wire \bit_sel_reg[59] ;
 wire \bit_sel_reg[5] ;
 wire \bit_sel_reg[60] ;
 wire \bit_sel_reg[61] ;
 wire \bit_sel_reg[62] ;
 wire \bit_sel_reg[63] ;
 wire \bit_sel_reg[6] ;
 wire \bit_sel_reg[7] ;
 wire \bit_sel_reg[8] ;
 wire \bit_sel_reg[9] ;
 wire \col_prog_n[0] ;
 wire \col_prog_n[10] ;
 wire \col_prog_n[11] ;
 wire \col_prog_n[12] ;
 wire \col_prog_n[13] ;
 wire \col_prog_n[14] ;
 wire \col_prog_n[15] ;
 wire \col_prog_n[1] ;
 wire \col_prog_n[2] ;
 wire \col_prog_n[3] ;
 wire \col_prog_n[4] ;
 wire \col_prog_n[5] ;
 wire \col_prog_n[6] ;
 wire \col_prog_n[7] ;
 wire \col_prog_n[8] ;
 wire \col_prog_n[9] ;
 wire \col_prog_n_reg[0] ;
 wire \col_prog_n_reg[10] ;
 wire \col_prog_n_reg[11] ;
 wire \col_prog_n_reg[12] ;
 wire \col_prog_n_reg[13] ;
 wire \col_prog_n_reg[14] ;
 wire \col_prog_n_reg[15] ;
 wire \col_prog_n_reg[1] ;
 wire \col_prog_n_reg[2] ;
 wire \col_prog_n_reg[3] ;
 wire \col_prog_n_reg[4] ;
 wire \col_prog_n_reg[5] ;
 wire \col_prog_n_reg[6] ;
 wire \col_prog_n_reg[7] ;
 wire \col_prog_n_reg[8] ;
 wire \col_prog_n_reg[9] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \efuse_out[0] ;
 wire \efuse_out[10] ;
 wire \efuse_out[11] ;
 wire \efuse_out[12] ;
 wire \efuse_out[13] ;
 wire \efuse_out[14] ;
 wire \efuse_out[15] ;
 wire \efuse_out[1] ;
 wire \efuse_out[2] ;
 wire \efuse_out[3] ;
 wire \efuse_out[4] ;
 wire \efuse_out[5] ;
 wire \efuse_out[6] ;
 wire \efuse_out[7] ;
 wire \efuse_out[8] ;
 wire \efuse_out[9] ;
 wire one;
 wire \preset_n[0] ;
 wire \preset_n[1] ;
 wire \preset_n_reg[0] ;
 wire \preset_n_reg[1] ;
 wire \sense[0] ;
 wire \sense[1] ;
 wire \sense_del[0] ;
 wire \sense_del[1] ;
 wire \sense_reg[0] ;
 wire \sense_reg[1] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0449_ (.I(\preset_n_reg[1] ),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0450_ (.I(\preset_n_reg[0] ),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0451_ (.I(\state[3] ),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0452_ (.I(\counter[9] ),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0453_ (.I(\counter[8] ),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0454_ (.I(\counter[7] ),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0455_ (.I(\counter[6] ),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0456_ (.I(\counter[5] ),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0457_ (.I(\counter[4] ),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0458_ (.I(\counter[3] ),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0459_ (.I(\counter[2] ),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0460_ (.I(\counter[1] ),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0461_ (.I(net21),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0462_ (.I(net29),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0463_ (.I(\state[1] ),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0464_ (.I(net28),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0465_ (.I(net27),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0466_ (.I(net26),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0467_ (.I(net25),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0468_ (.I(net24),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0469_ (.I(net23),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0470_ (.I(net22),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0471_ (.I(\sense_reg[1] ),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0472_ (.I(\sense_reg[0] ),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0473_ (.I(\state[0] ),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0474_ (.I(net7),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0475_ (.I(net6),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0476_ (.I(net1),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0477_ (.I(net2),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0478_ (.I(net3),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0479_ (.I(net4),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0480_ (.I(net5),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0481_ (.I(net17),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0482_ (.A1(net8),
    .A2(net19),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0483_ (.A1(net8),
    .A2(net19),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0484_ (.A1(net21),
    .A2(_0237_),
    .A3(net20),
    .A4(_0246_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0485_ (.I(_0247_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0486_ (.A1(_0237_),
    .A2(\state[2] ),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0487_ (.A1(_0247_),
    .A2(_0248_),
    .B(_0238_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0488_ (.A1(_0237_),
    .A2(_0000_),
    .B(\state[2] ),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0489_ (.A1(_0213_),
    .A2(_0249_),
    .B(_0250_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0490_ (.A1(_0247_),
    .A2(_0248_),
    .B(net7),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0491_ (.A1(_0214_),
    .A2(_0251_),
    .B(_0250_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0492_ (.A1(\state[3] ),
    .A2(net7),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0493_ (.A1(net18),
    .A2(net16),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0494_ (.A1(\col_prog_n_reg[15] ),
    .A2(_0252_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0495_ (.A1(\counter[2] ),
    .A2(\counter[1] ),
    .A3(\counter[0] ),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0496_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .A4(\counter[0] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0497_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .A3(\counter[5] ),
    .A4(\counter[4] ),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0498_ (.A1(_0256_),
    .A2(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0499_ (.A1(_0217_),
    .A2(_0256_),
    .A3(_0257_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0500_ (.A1(_0215_),
    .A2(\counter[9] ),
    .A3(_0259_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0501_ (.A1(\counter[9] ),
    .A2(\counter[8] ),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0502_ (.A1(\state[3] ),
    .A2(_0256_),
    .A3(_0257_),
    .A4(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0503_ (.A1(\state[3] ),
    .A2(_0256_),
    .A3(_0257_),
    .A4(_0261_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0504_ (.A1(_0252_),
    .A2(_0253_),
    .B(_0254_),
    .C(_0263_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0505_ (.A1(\col_prog_n_reg[14] ),
    .A2(_0252_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0506_ (.A1(net18),
    .A2(net15),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0507_ (.A1(_0252_),
    .A2(_0265_),
    .B(_0264_),
    .C(_0263_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0508_ (.A1(net18),
    .A2(net14),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0509_ (.A1(\col_prog_n_reg[13] ),
    .A2(_0252_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0510_ (.A1(_0252_),
    .A2(_0266_),
    .B(_0267_),
    .C(_0263_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0511_ (.A1(\col_prog_n_reg[12] ),
    .A2(_0252_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0512_ (.A1(net18),
    .A2(net13),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0513_ (.A1(_0252_),
    .A2(_0269_),
    .B(_0268_),
    .C(_0263_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0514_ (.A1(net18),
    .A2(net12),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0515_ (.A1(\col_prog_n_reg[11] ),
    .A2(_0252_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0516_ (.A1(_0252_),
    .A2(_0270_),
    .B(_0271_),
    .C(_0263_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0517_ (.A1(net18),
    .A2(net11),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0518_ (.A1(\col_prog_n_reg[10] ),
    .A2(_0252_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0519_ (.A1(_0252_),
    .A2(_0272_),
    .B(_0273_),
    .C(_0263_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0520_ (.A1(\col_prog_n_reg[9] ),
    .A2(_0252_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0521_ (.A1(net18),
    .A2(net10),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0522_ (.A1(_0252_),
    .A2(_0275_),
    .B(_0274_),
    .C(_0263_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0523_ (.A1(\col_prog_n_reg[8] ),
    .A2(_0252_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0524_ (.A1(net18),
    .A2(net9),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0525_ (.A1(_0252_),
    .A2(_0277_),
    .B(_0276_),
    .C(_0263_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0526_ (.A1(\state[3] ),
    .A2(_0238_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0527_ (.A1(\col_prog_n_reg[7] ),
    .A2(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0528_ (.A1(_0253_),
    .A2(_0278_),
    .B(_0279_),
    .C(_0260_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0529_ (.A1(\col_prog_n_reg[6] ),
    .A2(_0278_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0530_ (.A1(_0265_),
    .A2(_0278_),
    .B(_0280_),
    .C(_0260_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0531_ (.A1(\col_prog_n_reg[5] ),
    .A2(_0278_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0532_ (.A1(_0266_),
    .A2(_0278_),
    .B(_0281_),
    .C(_0260_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0533_ (.A1(\col_prog_n_reg[4] ),
    .A2(_0278_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0534_ (.A1(_0269_),
    .A2(_0278_),
    .B(_0282_),
    .C(_0260_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0535_ (.A1(\col_prog_n_reg[3] ),
    .A2(_0278_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0536_ (.A1(_0270_),
    .A2(_0278_),
    .B(_0283_),
    .C(_0260_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0537_ (.A1(\col_prog_n_reg[2] ),
    .A2(_0278_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0538_ (.A1(_0272_),
    .A2(_0278_),
    .B(_0284_),
    .C(_0260_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0539_ (.A1(\col_prog_n_reg[1] ),
    .A2(_0278_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0540_ (.A1(_0275_),
    .A2(_0278_),
    .B(_0285_),
    .C(_0260_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0541_ (.A1(\col_prog_n_reg[0] ),
    .A2(_0278_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0542_ (.A1(_0277_),
    .A2(_0278_),
    .B(_0286_),
    .C(_0260_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0543_ (.A1(\state[0] ),
    .A2(\state[2] ),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0544_ (.A1(\bit_sel_reg[63] ),
    .A2(net35),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0545_ (.A1(net1),
    .A2(net2),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0546_ (.A1(_0242_),
    .A2(_0243_),
    .A3(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0547_ (.A1(net5),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0548_ (.A1(_0225_),
    .A2(\state[0] ),
    .A3(net20),
    .A4(_0245_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0549_ (.A1(_0225_),
    .A2(\state[0] ),
    .A3(net20),
    .A4(_0245_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0550_ (.A1(\state[2] ),
    .A2(_0292_),
    .B(net6),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0551_ (.A1(_0291_),
    .A2(net32),
    .B(_0288_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0552_ (.A1(\bit_sel_reg[62] ),
    .A2(net36),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0553_ (.A1(net1),
    .A2(_0241_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0554_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0555_ (.A1(net34),
    .A2(_0297_),
    .B(_0295_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0556_ (.A1(\bit_sel_reg[61] ),
    .A2(net35),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0557_ (.A1(_0240_),
    .A2(net2),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0558_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0559_ (.A1(_0294_),
    .A2(_0300_),
    .B(_0298_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0560_ (.A1(\bit_sel_reg[60] ),
    .A2(net36),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0561_ (.A1(net1),
    .A2(net2),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0562_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0563_ (.A1(net34),
    .A2(_0303_),
    .B(_0301_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0564_ (.A1(\bit_sel_reg[59] ),
    .A2(net35),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0565_ (.A1(net3),
    .A2(_0289_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0566_ (.A1(net4),
    .A2(net5),
    .A3(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0567_ (.A1(net32),
    .A2(_0306_),
    .B(_0304_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0568_ (.A1(\bit_sel_reg[58] ),
    .A2(net35),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0569_ (.A1(net1),
    .A2(_0241_),
    .A3(net3),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0570_ (.A1(net4),
    .A2(net5),
    .A3(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0571_ (.A1(net34),
    .A2(_0309_),
    .B(_0307_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0572_ (.A1(\bit_sel_reg[57] ),
    .A2(_0287_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0573_ (.A1(_0240_),
    .A2(net2),
    .A3(net3),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0574_ (.A1(net4),
    .A2(net5),
    .A3(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0575_ (.A1(_0294_),
    .A2(_0312_),
    .B(_0310_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0576_ (.A1(\bit_sel_reg[56] ),
    .A2(net35),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0577_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0578_ (.A1(net4),
    .A2(net5),
    .A3(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0579_ (.A1(net33),
    .A2(_0315_),
    .B(_0313_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0580_ (.A1(\bit_sel_reg[55] ),
    .A2(net36),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0581_ (.A1(_0242_),
    .A2(net4),
    .A3(_0289_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0582_ (.A1(net5),
    .A2(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0583_ (.A1(net32),
    .A2(_0318_),
    .B(_0316_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0584_ (.A1(\bit_sel_reg[54] ),
    .A2(net36),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0585_ (.A1(net1),
    .A2(_0241_),
    .A3(_0242_),
    .A4(net4),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0586_ (.A1(net5),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0587_ (.A1(net34),
    .A2(_0321_),
    .B(_0319_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0588_ (.A1(\bit_sel_reg[53] ),
    .A2(_0287_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0589_ (.A1(_0240_),
    .A2(net2),
    .A3(_0242_),
    .A4(net4),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0590_ (.A1(net5),
    .A2(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0591_ (.A1(net33),
    .A2(_0324_),
    .B(_0322_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0592_ (.A1(\bit_sel_reg[52] ),
    .A2(net36),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0593_ (.A1(net3),
    .A2(_0243_),
    .A3(net5),
    .A4(_0302_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0594_ (.A1(net34),
    .A2(_0326_),
    .B(_0325_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0595_ (.A1(\bit_sel_reg[51] ),
    .A2(net35),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0596_ (.A1(net3),
    .A2(net4),
    .A3(_0289_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0597_ (.A1(net5),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0598_ (.A1(net33),
    .A2(_0329_),
    .B(_0327_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0599_ (.A1(\bit_sel_reg[50] ),
    .A2(net36),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0600_ (.A1(net1),
    .A2(_0241_),
    .A3(net3),
    .A4(net4),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0601_ (.A1(net5),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0602_ (.A1(net34),
    .A2(_0332_),
    .B(_0330_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0603_ (.A1(\bit_sel_reg[49] ),
    .A2(net35),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0604_ (.A1(_0240_),
    .A2(net2),
    .A3(net3),
    .A4(net4),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0605_ (.A1(net5),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0606_ (.A1(net33),
    .A2(_0335_),
    .B(_0333_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0607_ (.A1(\bit_sel_reg[48] ),
    .A2(net35),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0608_ (.A1(_0243_),
    .A2(_0314_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0609_ (.A1(net5),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0610_ (.A1(net33),
    .A2(_0338_),
    .B(_0336_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0611_ (.A1(\bit_sel_reg[47] ),
    .A2(net35),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0612_ (.A1(_0244_),
    .A2(_0290_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0613_ (.A1(net32),
    .A2(_0340_),
    .B(_0339_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0614_ (.A1(\bit_sel_reg[46] ),
    .A2(net36),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0615_ (.A1(net3),
    .A2(net4),
    .A3(_0244_),
    .A4(_0296_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0616_ (.A1(net34),
    .A2(_0342_),
    .B(_0341_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0617_ (.A1(\bit_sel_reg[45] ),
    .A2(net35),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0618_ (.A1(net3),
    .A2(net4),
    .A3(_0244_),
    .A4(_0299_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0619_ (.A1(_0294_),
    .A2(_0344_),
    .B(_0343_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0620_ (.A1(\bit_sel_reg[44] ),
    .A2(net35),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0621_ (.A1(net3),
    .A2(net4),
    .A3(_0244_),
    .A4(_0302_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0622_ (.A1(net32),
    .A2(_0346_),
    .B(_0345_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0623_ (.A1(\bit_sel_reg[43] ),
    .A2(net35),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0624_ (.A1(net4),
    .A2(_0244_),
    .A3(_0305_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0625_ (.A1(net32),
    .A2(_0348_),
    .B(_0347_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0626_ (.A1(\bit_sel_reg[42] ),
    .A2(net36),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0627_ (.A1(net4),
    .A2(_0244_),
    .A3(_0308_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0628_ (.A1(net34),
    .A2(_0350_),
    .B(_0349_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0629_ (.A1(\bit_sel_reg[41] ),
    .A2(_0287_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0630_ (.A1(net4),
    .A2(_0244_),
    .A3(_0311_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0631_ (.A1(_0294_),
    .A2(_0352_),
    .B(_0351_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0632_ (.A1(\bit_sel_reg[40] ),
    .A2(net35),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0633_ (.A1(net4),
    .A2(_0244_),
    .A3(_0314_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0634_ (.A1(net33),
    .A2(_0354_),
    .B(_0353_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0635_ (.A1(\bit_sel_reg[39] ),
    .A2(net36),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0636_ (.A1(_0244_),
    .A2(_0317_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0637_ (.A1(net32),
    .A2(_0356_),
    .B(_0355_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0638_ (.A1(\bit_sel_reg[38] ),
    .A2(net36),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0639_ (.A1(_0244_),
    .A2(_0320_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0640_ (.A1(net34),
    .A2(_0358_),
    .B(_0357_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0641_ (.A1(\bit_sel_reg[37] ),
    .A2(net35),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0642_ (.A1(_0244_),
    .A2(_0323_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0643_ (.A1(net33),
    .A2(_0360_),
    .B(_0359_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0644_ (.A1(\bit_sel_reg[36] ),
    .A2(net35),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0645_ (.A1(net3),
    .A2(_0243_),
    .A3(_0244_),
    .A4(_0302_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0646_ (.A1(net32),
    .A2(_0362_),
    .B(_0361_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0647_ (.A1(\bit_sel_reg[35] ),
    .A2(net35),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0648_ (.A1(_0244_),
    .A2(_0328_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0649_ (.A1(net33),
    .A2(_0364_),
    .B(_0363_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0650_ (.A1(\bit_sel_reg[34] ),
    .A2(net36),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0651_ (.A1(_0244_),
    .A2(_0331_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0652_ (.A1(net34),
    .A2(_0366_),
    .B(_0365_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0653_ (.A1(\bit_sel_reg[33] ),
    .A2(_0287_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0654_ (.A1(_0244_),
    .A2(_0334_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0655_ (.A1(net33),
    .A2(_0368_),
    .B(_0367_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0656_ (.A1(\bit_sel_reg[32] ),
    .A2(net35),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0657_ (.A1(_0244_),
    .A2(_0337_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0658_ (.A1(net33),
    .A2(_0370_),
    .B(_0369_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0659_ (.A1(\bit_sel_reg[31] ),
    .A2(net35),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0660_ (.A1(\state[2] ),
    .A2(_0292_),
    .B(_0239_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0661_ (.A1(_0291_),
    .A2(net30),
    .B(_0371_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0662_ (.A1(\bit_sel_reg[30] ),
    .A2(net36),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0663_ (.A1(_0297_),
    .A2(net31),
    .B(_0373_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0664_ (.A1(\bit_sel_reg[29] ),
    .A2(net36),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0665_ (.A1(_0300_),
    .A2(_0372_),
    .B(_0374_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0666_ (.A1(\bit_sel_reg[28] ),
    .A2(net36),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0667_ (.A1(_0303_),
    .A2(net31),
    .B(_0375_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0668_ (.A1(\bit_sel_reg[27] ),
    .A2(net35),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0669_ (.A1(_0306_),
    .A2(net30),
    .B(_0376_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0670_ (.A1(\bit_sel_reg[26] ),
    .A2(net35),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0671_ (.A1(_0309_),
    .A2(net30),
    .B(_0377_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0672_ (.A1(\bit_sel_reg[25] ),
    .A2(_0287_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0673_ (.A1(_0312_),
    .A2(_0372_),
    .B(_0378_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0674_ (.A1(\bit_sel_reg[24] ),
    .A2(net35),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0675_ (.A1(_0315_),
    .A2(_0372_),
    .B(_0379_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0676_ (.A1(\bit_sel_reg[23] ),
    .A2(net36),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0677_ (.A1(_0318_),
    .A2(net31),
    .B(_0380_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0678_ (.A1(\bit_sel_reg[22] ),
    .A2(net36),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0679_ (.A1(_0321_),
    .A2(net31),
    .B(_0381_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0680_ (.A1(\bit_sel_reg[21] ),
    .A2(_0287_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0681_ (.A1(_0324_),
    .A2(_0372_),
    .B(_0382_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0682_ (.A1(\bit_sel_reg[20] ),
    .A2(net36),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0683_ (.A1(_0326_),
    .A2(net31),
    .B(_0383_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0684_ (.A1(\bit_sel_reg[19] ),
    .A2(net35),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0685_ (.A1(_0329_),
    .A2(_0372_),
    .B(_0384_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0686_ (.A1(\bit_sel_reg[18] ),
    .A2(net36),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0687_ (.A1(_0332_),
    .A2(net31),
    .B(_0385_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0688_ (.A1(\bit_sel_reg[17] ),
    .A2(net35),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0689_ (.A1(_0335_),
    .A2(net30),
    .B(_0386_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0690_ (.A1(\bit_sel_reg[16] ),
    .A2(net35),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0691_ (.A1(_0338_),
    .A2(_0372_),
    .B(_0387_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0692_ (.A1(\bit_sel_reg[15] ),
    .A2(net35),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0693_ (.A1(_0340_),
    .A2(net30),
    .B(_0388_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0694_ (.A1(\bit_sel_reg[14] ),
    .A2(net36),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0695_ (.A1(_0342_),
    .A2(net30),
    .B(_0389_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0696_ (.A1(\bit_sel_reg[13] ),
    .A2(net36),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0697_ (.A1(_0344_),
    .A2(net31),
    .B(_0390_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0698_ (.A1(\bit_sel_reg[12] ),
    .A2(net35),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0699_ (.A1(_0346_),
    .A2(net30),
    .B(_0391_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0700_ (.A1(\bit_sel_reg[11] ),
    .A2(net35),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0701_ (.A1(_0348_),
    .A2(net30),
    .B(_0392_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0702_ (.A1(\bit_sel_reg[10] ),
    .A2(net36),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0703_ (.A1(_0350_),
    .A2(net31),
    .B(_0393_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0704_ (.A1(\bit_sel_reg[9] ),
    .A2(_0287_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0705_ (.A1(_0352_),
    .A2(_0372_),
    .B(_0394_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0706_ (.A1(\bit_sel_reg[8] ),
    .A2(net35),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0707_ (.A1(_0354_),
    .A2(_0372_),
    .B(_0395_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0708_ (.A1(\bit_sel_reg[7] ),
    .A2(net36),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0709_ (.A1(_0356_),
    .A2(net31),
    .B(_0396_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0710_ (.A1(\bit_sel_reg[6] ),
    .A2(net36),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0711_ (.A1(_0358_),
    .A2(net31),
    .B(_0397_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0712_ (.A1(\bit_sel_reg[5] ),
    .A2(net35),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0713_ (.A1(_0360_),
    .A2(_0372_),
    .B(_0398_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0714_ (.A1(\bit_sel_reg[4] ),
    .A2(net35),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0715_ (.A1(_0362_),
    .A2(net30),
    .B(_0399_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0716_ (.A1(\bit_sel_reg[3] ),
    .A2(net35),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0717_ (.A1(_0364_),
    .A2(_0372_),
    .B(_0400_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0718_ (.A1(\bit_sel_reg[2] ),
    .A2(net36),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0719_ (.A1(_0366_),
    .A2(net31),
    .B(_0401_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0720_ (.A1(\bit_sel_reg[1] ),
    .A2(_0287_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0721_ (.A1(_0368_),
    .A2(_0372_),
    .B(_0402_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0722_ (.A1(\bit_sel_reg[0] ),
    .A2(net35),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0723_ (.A1(_0370_),
    .A2(_0372_),
    .B(_0403_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0724_ (.A1(_0215_),
    .A2(\state[0] ),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0725_ (.A1(\state[3] ),
    .A2(_0237_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0726_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0259_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0727_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0262_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0728_ (.A1(_0292_),
    .A2(_0404_),
    .B(_0263_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0729_ (.A1(_0215_),
    .A2(_0292_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0730_ (.A1(_0216_),
    .A2(_0406_),
    .B(_0409_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0731_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0258_),
    .C(_0262_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0732_ (.A1(\state[3] ),
    .A2(_0259_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0733_ (.A1(_0217_),
    .A2(_0410_),
    .B1(_0411_),
    .B2(_0408_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0734_ (.A1(\state[0] ),
    .A2(_0293_),
    .B(_0262_),
    .C(_0215_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0735_ (.A1(_0237_),
    .A2(_0292_),
    .B(_0263_),
    .C(\state[3] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0736_ (.A1(_0221_),
    .A2(_0256_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0737_ (.A1(_0220_),
    .A2(_0221_),
    .A3(_0256_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0738_ (.A1(_0219_),
    .A2(_0220_),
    .A3(_0221_),
    .A4(_0256_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0739_ (.A1(\counter[7] ),
    .A2(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0740_ (.A1(_0292_),
    .A2(_0404_),
    .B1(_0416_),
    .B2(_0215_),
    .C(_0263_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0741_ (.A1(_0412_),
    .A2(_0417_),
    .B1(_0418_),
    .B2(_0218_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0742_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0415_),
    .C(_0262_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0743_ (.A1(_0219_),
    .A2(_0419_),
    .B(_0418_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0744_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0414_),
    .C(_0262_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0745_ (.A1(_0408_),
    .A2(_0415_),
    .B1(_0420_),
    .B2(_0220_),
    .C(_0409_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0746_ (.A1(_0215_),
    .A2(_0256_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0747_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0421_),
    .C(_0262_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0748_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0422_),
    .B2(_0221_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0749_ (.A1(_0293_),
    .A2(_0405_),
    .B(_0255_),
    .C(_0262_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0750_ (.A1(_0408_),
    .A2(_0421_),
    .B1(_0423_),
    .B2(_0222_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0751_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .B(\counter[2] ),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0752_ (.A1(_0255_),
    .A2(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0753_ (.A1(_0223_),
    .A2(_0407_),
    .B1(_0413_),
    .B2(_0425_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0754_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0755_ (.A1(_0224_),
    .A2(_0407_),
    .B1(_0413_),
    .B2(_0426_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0756_ (.I0(_0412_),
    .I1(_0408_),
    .S(\counter[0] ),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0757_ (.A1(\state[3] ),
    .A2(_0263_),
    .B(_0237_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0758_ (.A1(\state[3] ),
    .A2(_0227_),
    .B1(_0427_),
    .B2(_0225_),
    .C(_0260_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0759_ (.A1(net7),
    .A2(\efuse_out[15] ),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0760_ (.A1(_0238_),
    .A2(\efuse_out[7] ),
    .B(_0227_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0761_ (.A1(_0226_),
    .A2(_0227_),
    .B1(_0428_),
    .B2(_0429_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0762_ (.A1(net7),
    .A2(\efuse_out[14] ),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0763_ (.A1(_0238_),
    .A2(\efuse_out[6] ),
    .B(_0227_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0764_ (.A1(_0227_),
    .A2(_0228_),
    .B1(_0430_),
    .B2(_0431_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0765_ (.A1(net7),
    .A2(\efuse_out[13] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0766_ (.A1(_0238_),
    .A2(\efuse_out[5] ),
    .B(_0227_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0767_ (.A1(_0227_),
    .A2(_0229_),
    .B1(_0432_),
    .B2(_0433_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0768_ (.A1(net7),
    .A2(\efuse_out[12] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0769_ (.A1(_0238_),
    .A2(\efuse_out[4] ),
    .B(_0227_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0770_ (.A1(_0227_),
    .A2(_0230_),
    .B1(_0434_),
    .B2(_0435_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0771_ (.A1(net7),
    .A2(\efuse_out[11] ),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0772_ (.A1(_0238_),
    .A2(\efuse_out[3] ),
    .B(_0227_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0773_ (.A1(_0227_),
    .A2(_0231_),
    .B1(_0436_),
    .B2(_0437_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0774_ (.A1(net7),
    .A2(\efuse_out[10] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0775_ (.A1(_0238_),
    .A2(\efuse_out[2] ),
    .B(_0227_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0776_ (.A1(_0227_),
    .A2(_0232_),
    .B1(_0438_),
    .B2(_0439_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0777_ (.A1(net7),
    .A2(\efuse_out[9] ),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0778_ (.A1(_0238_),
    .A2(\efuse_out[1] ),
    .B(_0227_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0779_ (.A1(_0227_),
    .A2(_0233_),
    .B1(_0440_),
    .B2(_0441_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0780_ (.A1(net7),
    .A2(\efuse_out[8] ),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0781_ (.A1(_0238_),
    .A2(\efuse_out[0] ),
    .B(_0227_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0782_ (.A1(_0227_),
    .A2(_0234_),
    .B1(_0442_),
    .B2(_0443_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0783_ (.A1(_0227_),
    .A2(\state[0] ),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0784_ (.A1(_0000_),
    .A2(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0785_ (.A1(_0000_),
    .A2(_0444_),
    .B(net7),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0786_ (.A1(\state[1] ),
    .A2(_0445_),
    .B1(_0446_),
    .B2(_0235_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0787_ (.A1(_0000_),
    .A2(_0444_),
    .B(_0238_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0788_ (.A1(\state[1] ),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0236_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0789_ (.A1(net21),
    .A2(_0246_),
    .B(\state[0] ),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0790_ (.A1(_0227_),
    .A2(_0263_),
    .A3(_0448_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0791_ (.A1(_0215_),
    .A2(_0262_),
    .B(_0293_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0792_ (.I(net37),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0793_ (.I(net37),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0794_ (.I(net38),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0795_ (.I(net37),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0796_ (.I(net38),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0797_ (.I(net37),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0798_ (.I(net38),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0799_ (.I(net38),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0800_ (.I(net38),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0801_ (.I(net38),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0802_ (.I(net38),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0803_ (.I(net38),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0804_ (.I(net17),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0805_ (.I(net17),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0806_ (.I(net17),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0807_ (.I(net17),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0808_ (.I(net17),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0809_ (.I(net17),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0810_ (.I(net38),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0811_ (.I(net38),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0812_ (.I(net38),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0813_ (.I(net38),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0814_ (.I(net17),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0815_ (.I(net38),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0816_ (.I(net38),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0817_ (.I(net38),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0818_ (.I(net37),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0819_ (.I(net38),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0820_ (.I(net37),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0821_ (.I(net37),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0822_ (.I(net37),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0823_ (.I(net37),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0824_ (.I(net38),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0825_ (.I(net38),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0826_ (.I(net37),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0827_ (.I(net37),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0828_ (.I(net37),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0829_ (.I(net37),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0830_ (.I(net37),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0831_ (.I(net37),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0832_ (.I(net38),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0833_ (.I(net37),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0834_ (.I(net37),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0835_ (.I(net38),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0836_ (.I(net37),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0837_ (.I(net38),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0838_ (.I(net37),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0839_ (.I(net37),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0840_ (.I(net38),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0841_ (.I(net38),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0842_ (.I(net37),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0843_ (.I(net37),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0844_ (.I(net37),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0845_ (.I(net37),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0846_ (.I(net37),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0847_ (.I(net37),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0848_ (.I(net38),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0849_ (.I(net38),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0850_ (.I(net37),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0851_ (.I(net38),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0852_ (.I(net37),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0853_ (.I(net37),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0854_ (.I(net37),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0855_ (.I(net37),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0856_ (.I(net38),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0857_ (.I(net38),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0858_ (.I(net37),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0859_ (.I(net37),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0860_ (.I(net37),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0861_ (.I(net37),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0862_ (.I(net37),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0863_ (.I(net37),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0864_ (.I(net38),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0865_ (.I(net37),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0866_ (.I(net37),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0867_ (.I(net38),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0868_ (.I(net37),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0869_ (.I(net38),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0870_ (.I(net37),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0871_ (.I(net37),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0872_ (.I(net38),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0873_ (.I(net38),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0874_ (.I(net37),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0875_ (.I(net37),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0876_ (.I(net37),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0877_ (.I(net37),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0878_ (.I(net37),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0879_ (.I(net37),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0880_ (.I(net37),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0881_ (.I(net37),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0882_ (.I(net37),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0883_ (.I(net38),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0884_ (.I(net38),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0885_ (.I(net38),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0886_ (.I(net37),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0887_ (.I(net38),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0888_ (.I(net38),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0889_ (.I(net38),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0890_ (.I(net17),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0891_ (.I(net17),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0892_ (.I(net38),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0893_ (.I(net38),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0894_ (.I(net17),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0895_ (.I(net17),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0896_ (.I(net37),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0897_ (.I(net38),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0898_ (.D(_0001_),
    .SETN(_0003_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0899_ (.D(\state[2] ),
    .RN(_0004_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0900_ (.D(_0000_),
    .RN(_0005_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0901_ (.D(_0002_),
    .RN(_0006_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0902_ (.D(_0110_),
    .RN(_0007_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\sense_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0903_ (.D(_0111_),
    .RN(_0008_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\sense_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0904_ (.D(_0112_),
    .RN(_0009_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0905_ (.D(_0113_),
    .RN(_0010_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0906_ (.D(_0114_),
    .RN(_0011_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0907_ (.D(_0115_),
    .RN(_0012_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0908_ (.D(_0116_),
    .RN(_0013_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0909_ (.D(_0117_),
    .RN(_0014_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0910_ (.D(_0118_),
    .RN(_0015_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0911_ (.D(_0119_),
    .RN(_0016_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0912_ (.D(_0120_),
    .RN(_0017_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0913_ (.D(_0121_),
    .RN(_0018_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0914_ (.D(_0122_),
    .RN(_0019_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0915_ (.D(_0123_),
    .RN(_0020_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0916_ (.D(_0124_),
    .RN(_0021_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0917_ (.D(_0125_),
    .RN(_0022_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0918_ (.D(_0126_),
    .RN(_0023_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0919_ (.D(_0127_),
    .RN(_0024_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0920_ (.D(_0128_),
    .RN(_0025_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0921_ (.D(_0129_),
    .RN(_0026_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0922_ (.D(_0130_),
    .RN(_0027_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0923_ (.D(_0131_),
    .RN(_0028_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0924_ (.D(_0132_),
    .RN(_0029_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0925_ (.D(_0133_),
    .RN(_0030_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0926_ (.D(_0134_),
    .RN(_0031_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0927_ (.D(_0135_),
    .RN(_0032_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0928_ (.D(_0136_),
    .RN(_0033_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0929_ (.D(_0137_),
    .RN(_0034_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0930_ (.D(_0138_),
    .RN(_0035_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0931_ (.D(_0139_),
    .RN(_0036_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0932_ (.D(_0140_),
    .RN(_0037_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0933_ (.D(_0141_),
    .RN(_0038_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0934_ (.D(_0142_),
    .RN(_0039_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0935_ (.D(_0143_),
    .RN(_0040_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0936_ (.D(_0144_),
    .RN(_0041_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0937_ (.D(_0145_),
    .RN(_0042_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0938_ (.D(_0146_),
    .RN(_0043_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0939_ (.D(_0147_),
    .RN(_0044_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0940_ (.D(_0148_),
    .RN(_0045_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0941_ (.D(_0149_),
    .RN(_0046_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0942_ (.D(_0150_),
    .RN(_0047_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0943_ (.D(_0151_),
    .RN(_0048_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0944_ (.D(_0152_),
    .RN(_0049_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0945_ (.D(_0153_),
    .RN(_0050_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0946_ (.D(_0154_),
    .RN(_0051_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0947_ (.D(_0155_),
    .RN(_0052_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0948_ (.D(_0156_),
    .RN(_0053_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0949_ (.D(_0157_),
    .RN(_0054_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0950_ (.D(_0158_),
    .RN(_0055_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0951_ (.D(_0159_),
    .RN(_0056_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0952_ (.D(_0160_),
    .RN(_0057_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0953_ (.D(_0161_),
    .RN(_0058_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0954_ (.D(_0162_),
    .RN(_0059_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0955_ (.D(_0163_),
    .RN(_0060_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0956_ (.D(_0164_),
    .RN(_0061_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0957_ (.D(_0165_),
    .RN(_0062_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0958_ (.D(_0166_),
    .RN(_0063_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0959_ (.D(_0167_),
    .RN(_0064_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0960_ (.D(_0168_),
    .RN(_0065_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0961_ (.D(_0169_),
    .RN(_0066_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0962_ (.D(_0170_),
    .RN(_0067_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0963_ (.D(_0171_),
    .RN(_0068_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0964_ (.D(_0172_),
    .RN(_0069_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0965_ (.D(_0173_),
    .RN(_0070_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0966_ (.D(_0174_),
    .RN(_0071_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0967_ (.D(_0175_),
    .RN(_0072_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0968_ (.D(_0176_),
    .RN(_0073_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0969_ (.D(_0177_),
    .RN(_0074_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0970_ (.D(_0178_),
    .RN(_0075_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0971_ (.D(_0179_),
    .RN(_0076_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0972_ (.D(_0180_),
    .RN(_0077_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0973_ (.D(_0181_),
    .RN(_0078_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0974_ (.D(_0182_),
    .RN(_0079_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0975_ (.D(_0183_),
    .RN(_0080_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0976_ (.D(_0184_),
    .RN(_0081_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0977_ (.D(_0185_),
    .RN(_0082_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0978_ (.D(_0186_),
    .RN(_0083_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\bit_sel_reg[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0979_ (.D(_0187_),
    .RN(_0084_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0980_ (.D(_0188_),
    .RN(_0085_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\bit_sel_reg[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0981_ (.D(_0189_),
    .RN(_0086_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0982_ (.D(_0190_),
    .RN(_0087_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0983_ (.D(_0191_),
    .RN(_0088_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0984_ (.D(_0192_),
    .RN(_0089_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0985_ (.D(_0193_),
    .RN(_0090_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\bit_sel_reg[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _0986_ (.D(_0194_),
    .RN(_0091_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\bit_sel_reg[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0987_ (.D(_0195_),
    .SETN(_0092_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0988_ (.D(_0196_),
    .SETN(_0093_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0989_ (.D(_0197_),
    .SETN(_0094_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0990_ (.D(_0198_),
    .SETN(_0095_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0991_ (.D(_0199_),
    .SETN(_0096_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0992_ (.D(_0200_),
    .SETN(_0097_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0993_ (.D(_0201_),
    .SETN(_0098_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0994_ (.D(_0202_),
    .SETN(_0099_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0995_ (.D(_0203_),
    .SETN(_0100_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0996_ (.D(_0204_),
    .SETN(_0101_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0997_ (.D(_0205_),
    .SETN(_0102_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0998_ (.D(_0206_),
    .SETN(_0103_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _0999_ (.D(_0207_),
    .SETN(_0104_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1000_ (.D(_0208_),
    .SETN(_0105_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1001_ (.D(_0209_),
    .SETN(_0106_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1002_ (.D(_0210_),
    .SETN(_0107_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\col_prog_n_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1003_ (.D(_0211_),
    .SETN(_0108_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\preset_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1004_ (.D(_0212_),
    .SETN(_0109_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\preset_n_reg[1] ));
 efuse_array_64x8 \efuse_gen_depth[0].efuse_array  (.PRESET_N(\preset_n[0] ),
    .SENSE(\sense[0] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[7] ,
    \col_prog_n[6] ,
    \col_prog_n[5] ,
    \col_prog_n[4] ,
    \col_prog_n[3] ,
    \col_prog_n[2] ,
    \col_prog_n[1] ,
    \col_prog_n[0] }),
    .OUT({\efuse_out[7] ,
    \efuse_out[6] ,
    \efuse_out[5] ,
    \efuse_out[4] ,
    \efuse_out[3] ,
    \efuse_out[2] ,
    \efuse_out[1] ,
    \efuse_out[0] }));
 efuse_array_64x8 \efuse_gen_depth[1].efuse_array  (.PRESET_N(\preset_n[1] ),
    .SENSE(\sense[1] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[15] ,
    \col_prog_n[14] ,
    \col_prog_n[13] ,
    \col_prog_n[12] ,
    \col_prog_n[11] ,
    \col_prog_n[10] ,
    \col_prog_n[9] ,
    \col_prog_n[8] }),
    .OUT({\efuse_out[15] ,
    \efuse_out[14] ,
    \efuse_out[13] ,
    \efuse_out[12] ,
    \efuse_out[11] ,
    \efuse_out[10] ,
    \efuse_out[9] ,
    \efuse_out[8] }));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[0].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[0] ),
    .S(write_enable_i),
    .Z(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[10].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[10] ),
    .S(write_enable_i),
    .Z(\col_prog_n[10] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[11].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[11] ),
    .S(write_enable_i),
    .Z(\col_prog_n[11] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[12].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[12] ),
    .S(write_enable_i),
    .Z(\col_prog_n[12] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[13].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[13] ),
    .S(write_enable_i),
    .Z(\col_prog_n[13] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[14].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[14] ),
    .S(write_enable_i),
    .Z(\col_prog_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[15].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[15] ),
    .S(write_enable_i),
    .Z(\col_prog_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[1].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[1] ),
    .S(write_enable_i),
    .Z(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[2].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[2] ),
    .S(write_enable_i),
    .Z(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[3].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[3] ),
    .S(write_enable_i),
    .Z(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[4].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[4] ),
    .S(write_enable_i),
    .Z(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[5].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[5] ),
    .S(write_enable_i),
    .Z(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[6].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[6] ),
    .S(write_enable_i),
    .Z(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[7].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[7] ),
    .S(write_enable_i),
    .Z(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[8].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[8] ),
    .S(write_enable_i),
    .Z(\col_prog_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[9].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[9] ),
    .S(write_enable_i),
    .Z(\col_prog_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[0].bitsel_buf_keep_cell  (.I(\bit_sel_reg[0] ),
    .Z(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[10].bitsel_buf_keep_cell  (.I(\bit_sel_reg[10] ),
    .Z(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[11].bitsel_buf_keep_cell  (.I(\bit_sel_reg[11] ),
    .Z(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[12].bitsel_buf_keep_cell  (.I(\bit_sel_reg[12] ),
    .Z(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[13].bitsel_buf_keep_cell  (.I(\bit_sel_reg[13] ),
    .Z(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[14].bitsel_buf_keep_cell  (.I(\bit_sel_reg[14] ),
    .Z(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[15].bitsel_buf_keep_cell  (.I(\bit_sel_reg[15] ),
    .Z(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[16].bitsel_buf_keep_cell  (.I(\bit_sel_reg[16] ),
    .Z(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[17].bitsel_buf_keep_cell  (.I(\bit_sel_reg[17] ),
    .Z(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[18].bitsel_buf_keep_cell  (.I(\bit_sel_reg[18] ),
    .Z(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[19].bitsel_buf_keep_cell  (.I(\bit_sel_reg[19] ),
    .Z(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[1].bitsel_buf_keep_cell  (.I(\bit_sel_reg[1] ),
    .Z(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[20].bitsel_buf_keep_cell  (.I(\bit_sel_reg[20] ),
    .Z(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[21].bitsel_buf_keep_cell  (.I(\bit_sel_reg[21] ),
    .Z(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[22].bitsel_buf_keep_cell  (.I(\bit_sel_reg[22] ),
    .Z(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[23].bitsel_buf_keep_cell  (.I(\bit_sel_reg[23] ),
    .Z(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[24].bitsel_buf_keep_cell  (.I(\bit_sel_reg[24] ),
    .Z(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[25].bitsel_buf_keep_cell  (.I(\bit_sel_reg[25] ),
    .Z(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[26].bitsel_buf_keep_cell  (.I(\bit_sel_reg[26] ),
    .Z(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[27].bitsel_buf_keep_cell  (.I(\bit_sel_reg[27] ),
    .Z(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[28].bitsel_buf_keep_cell  (.I(\bit_sel_reg[28] ),
    .Z(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[29].bitsel_buf_keep_cell  (.I(\bit_sel_reg[29] ),
    .Z(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[2].bitsel_buf_keep_cell  (.I(\bit_sel_reg[2] ),
    .Z(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[30].bitsel_buf_keep_cell  (.I(\bit_sel_reg[30] ),
    .Z(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[31].bitsel_buf_keep_cell  (.I(\bit_sel_reg[31] ),
    .Z(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[32].bitsel_buf_keep_cell  (.I(\bit_sel_reg[32] ),
    .Z(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[33].bitsel_buf_keep_cell  (.I(\bit_sel_reg[33] ),
    .Z(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[34].bitsel_buf_keep_cell  (.I(\bit_sel_reg[34] ),
    .Z(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[35].bitsel_buf_keep_cell  (.I(\bit_sel_reg[35] ),
    .Z(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[36].bitsel_buf_keep_cell  (.I(\bit_sel_reg[36] ),
    .Z(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[37].bitsel_buf_keep_cell  (.I(\bit_sel_reg[37] ),
    .Z(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[38].bitsel_buf_keep_cell  (.I(\bit_sel_reg[38] ),
    .Z(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[39].bitsel_buf_keep_cell  (.I(\bit_sel_reg[39] ),
    .Z(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[3].bitsel_buf_keep_cell  (.I(\bit_sel_reg[3] ),
    .Z(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[40].bitsel_buf_keep_cell  (.I(\bit_sel_reg[40] ),
    .Z(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[41].bitsel_buf_keep_cell  (.I(\bit_sel_reg[41] ),
    .Z(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[42].bitsel_buf_keep_cell  (.I(\bit_sel_reg[42] ),
    .Z(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[43].bitsel_buf_keep_cell  (.I(\bit_sel_reg[43] ),
    .Z(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[44].bitsel_buf_keep_cell  (.I(\bit_sel_reg[44] ),
    .Z(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[45].bitsel_buf_keep_cell  (.I(\bit_sel_reg[45] ),
    .Z(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[46].bitsel_buf_keep_cell  (.I(\bit_sel_reg[46] ),
    .Z(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[47].bitsel_buf_keep_cell  (.I(\bit_sel_reg[47] ),
    .Z(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[48].bitsel_buf_keep_cell  (.I(\bit_sel_reg[48] ),
    .Z(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[49].bitsel_buf_keep_cell  (.I(\bit_sel_reg[49] ),
    .Z(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[4].bitsel_buf_keep_cell  (.I(\bit_sel_reg[4] ),
    .Z(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[50].bitsel_buf_keep_cell  (.I(\bit_sel_reg[50] ),
    .Z(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[51].bitsel_buf_keep_cell  (.I(\bit_sel_reg[51] ),
    .Z(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[52].bitsel_buf_keep_cell  (.I(\bit_sel_reg[52] ),
    .Z(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[53].bitsel_buf_keep_cell  (.I(\bit_sel_reg[53] ),
    .Z(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[54].bitsel_buf_keep_cell  (.I(\bit_sel_reg[54] ),
    .Z(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[55].bitsel_buf_keep_cell  (.I(\bit_sel_reg[55] ),
    .Z(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[56].bitsel_buf_keep_cell  (.I(\bit_sel_reg[56] ),
    .Z(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[57].bitsel_buf_keep_cell  (.I(\bit_sel_reg[57] ),
    .Z(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[58].bitsel_buf_keep_cell  (.I(\bit_sel_reg[58] ),
    .Z(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[59].bitsel_buf_keep_cell  (.I(\bit_sel_reg[59] ),
    .Z(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[5].bitsel_buf_keep_cell  (.I(\bit_sel_reg[5] ),
    .Z(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[60].bitsel_buf_keep_cell  (.I(\bit_sel_reg[60] ),
    .Z(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[61].bitsel_buf_keep_cell  (.I(\bit_sel_reg[61] ),
    .Z(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[62].bitsel_buf_keep_cell  (.I(\bit_sel_reg[62] ),
    .Z(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[63].bitsel_buf_keep_cell  (.I(\bit_sel_reg[63] ),
    .Z(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[6].bitsel_buf_keep_cell  (.I(\bit_sel_reg[6] ),
    .Z(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[7].bitsel_buf_keep_cell  (.I(\bit_sel_reg[7] ),
    .Z(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[8].bitsel_buf_keep_cell  (.I(\bit_sel_reg[8] ),
    .Z(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[9].bitsel_buf_keep_cell  (.I(\bit_sel_reg[9] ),
    .Z(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].preset_buf_keep_cell  (.I(\preset_n_reg[0] ),
    .Z(\preset_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].sense_buf_keep_cell  (.I(\sense_del[0] ),
    .Z(\sense[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[0].sense_dly_keep_cell  (.I(\sense_reg[0] ),
    .Z(\sense_del[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[1].preset_buf_keep_cell  (.I(\preset_n_reg[1] ),
    .Z(\preset_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[1].sense_buf_keep_cell  (.I(\sense_del[1] ),
    .Z(\sense[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[1].sense_dly_keep_cell  (.I(\sense_reg[1] ),
    .Z(\sense_del[1] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh tie_keep_cell (.Z(one));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Left_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Left_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Left_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Left_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Left_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Left_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Left_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Left_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Left_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Left_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Left_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Left_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Left_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Left_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Left_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Left_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_3_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_3_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_3_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_3_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_3_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_3_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_3_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_3_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_3_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_3_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_3_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_3_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_3_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_3_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_3_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_3_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_3_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_3_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_3_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_3_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_3_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_3_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_3_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_3_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_3_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_3_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_3_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_3_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_3_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_3_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_3_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_3_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_3_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_3_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_3_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_3_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_3_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_3_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_3_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_3_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_3_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_3_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_3_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_3_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_3_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_3_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_3_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_3_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_3_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_3_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_3_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_3_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_3_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_3_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_3_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_3_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_3_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_3_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_3_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_3_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_3_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_3_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_3_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_3_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_3_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_3_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_3_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_3_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_3_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_3_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_3_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_3_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_3_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_3_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_3_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_3_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_3_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_3_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_3_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_3_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_3_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_3_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_3_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_3_Right_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_3_Right_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_3_Right_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_3_Right_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_3_Right_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_3_Right_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_3_Right_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_3_Right_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_3_Right_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_3_Right_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_3_Right_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_3_Right_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_3_Right_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_3_Right_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_3_Right_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_3_Right_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_3_Right_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_3_Right_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_3_Right_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_3_Right_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_3_Right_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_3_Right_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_3_Right_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_3_Right_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_3_Right_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_3_Right_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_3_Right_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_3_Right_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_3_Right_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_3_Right_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_3_Right_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_3_Right_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_3_Right_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_3_Right_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_3_Right_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_3_Right_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_3_Right_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_3_Right_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_3_Right_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_3_Right_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_3_Right_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_3_Right_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_3_Right_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_3_Right_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_3_Right_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_3_Right_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_3_Right_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_3_Right_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_3_Right_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_3_Right_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_3_Right_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_3_Right_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_3_Right_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_3_Right_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_3_Right_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_3_Right_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_3_Right_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_3_Right_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_3_Right_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_3_Right_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_3_Right_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_3_Right_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_3_Right_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_3_Right_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_3_Right_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_3_Right_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_3_Right_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_3_Right_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_3_Right_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_3_Right_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_3_Right_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_3_Right_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_3_Right_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_3_Right_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_3_Right_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_3_Right_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_3_Right_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_3_Right_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_3_Right_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_3_Right_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_3_Right_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_3_Right_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_3_Right_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_2_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_3_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_3_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_3_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_3_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_3_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_3_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_3_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_3_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_3_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_3_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_3_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_3_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_3_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_3_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_3_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_3_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_3_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_3_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_3_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_3_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_3_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_3_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_3_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_3_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_3_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_3_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_3_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_3_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_3_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_3_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_3_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_3_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_3_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_3_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_3_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_3_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_3_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_3_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_3_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_3_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_3_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_3_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_3_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_3_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_3_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_3_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_3_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_3_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_3_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_3_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_3_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_3_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_3_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_3_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_3_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_3_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_3_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_3_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_3_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_3_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_3_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_3_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_3_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_3_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_3_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_3_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_3_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_3_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_3_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_3_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_3_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_3_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_3_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_3_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_3_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_3_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_3_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_3_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_3_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_3_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_3_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_3_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_3_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_3_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_3_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_3_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_3_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_3_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_3_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_3_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_3_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_3_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_3_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_3_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_3_660 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(wb_adr_i[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(wb_adr_i[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(wb_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(wb_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(wb_adr_i[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(wb_adr_i[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(wb_adr_i[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(wb_cyc_i),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(wb_dat_i[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(wb_dat_i[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(wb_dat_i[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(wb_dat_i[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(wb_dat_i[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(wb_dat_i[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(wb_dat_i[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(wb_dat_i[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(wb_rst_i),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(wb_sel_i),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(wb_stb_i),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(wb_we_i),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output21 (.I(net21),
    .Z(wb_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output22 (.I(net22),
    .Z(wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output23 (.I(net23),
    .Z(wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output24 (.I(net24),
    .Z(wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output25 (.I(net25),
    .Z(wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output26 (.I(net26),
    .Z(wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output27 (.I(net27),
    .Z(wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output28 (.I(net28),
    .Z(wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output29 (.I(net29),
    .Z(wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap31 (.I(_0372_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap32 (.I(net34),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap34 (.I(_0294_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap35 (.I(_0287_),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap36 (.I(_0287_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew38 (.I(net17),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload0 (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload1 (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload2 (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 clkload3 (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload4 (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 clkload5 (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload6 (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_790 ();
endmodule
