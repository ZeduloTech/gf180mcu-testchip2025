VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180_ram_512x8_wrapper
  CLASS BLOCK ;
  FOREIGN gf180_ram_512x8_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 431.860 BY 484.880 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.215 0.000 172.335 29.595 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.760 0.000 163.880 29.595 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.295 0.000 155.415 29.595 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 281.325 0.000 282.445 18.645 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 275.820 0.000 276.940 12.700 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 272.085 0.000 273.205 15.120 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 268.860 0.000 269.980 17.355 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.525 0.000 149.645 15.020 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 145.030 0.000 146.150 12.620 ;
    END
  END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 251.710 0.000 252.830 36.390 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 44.706600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.680 0.000 140.800 16.615 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.320 0.000 10.440 25.675 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.030 0.000 62.150 8.505 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.270 0.000 68.390 8.505 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.975 0.000 120.095 16.910 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 307.235 0.000 308.355 25.675 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 358.910 0.000 360.030 8.505 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 365.150 0.000 366.270 8.505 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 416.860 0.000 417.980 25.675 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 14.466000 ;
    PORT
      LAYER Metal2 ;
        RECT 202.940 0.000 204.060 16.150 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.900 0.000 18.020 8.505 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.665 0.000 58.785 8.505 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.635 0.000 71.755 8.505 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.395 0.000 112.515 8.505 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 314.790 0.000 315.910 8.505 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 355.545 0.000 356.665 8.505 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 368.515 0.000 369.635 8.505 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 409.275 0.000 410.395 8.505 ;
    END
  END Q[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 0.000 2.000 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.800 0.000 428.800 482.160 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 3.000 0.000 5.000 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 429.800 0.000 431.800 482.160 ;
    END
  END VSS
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.695 0.000 13.815 8.185 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.020 0.000 64.140 8.185 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.270 0.000 66.390 8.185 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.020 0.000 118.140 8.185 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 310.575 0.000 311.695 8.185 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 360.900 0.000 362.020 8.185 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 363.150 0.000 364.270 8.185 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 413.475 0.000 414.595 8.185 ;
    END
  END WEN[7]
  OBS
      LAYER Nwell ;
        RECT 8.870 8.245 422.170 477.950 ;
      LAYER Metal1 ;
        RECT 1.410 1.410 430.450 483.470 ;
      LAYER Metal2 ;
        RECT 1.410 36.690 430.450 483.470 ;
        RECT 1.410 29.895 251.410 36.690 ;
        RECT 1.410 25.975 153.995 29.895 ;
        RECT 1.410 1.410 9.020 25.975 ;
        RECT 10.740 17.210 153.995 25.975 ;
        RECT 10.740 8.805 118.675 17.210 ;
        RECT 10.740 8.485 16.600 8.805 ;
        RECT 10.740 1.410 12.395 8.485 ;
        RECT 14.115 1.410 16.600 8.485 ;
        RECT 18.320 1.410 57.365 8.805 ;
        RECT 59.085 1.410 60.730 8.805 ;
        RECT 62.450 8.485 66.970 8.805 ;
        RECT 62.450 1.410 62.720 8.485 ;
        RECT 64.440 1.410 64.970 8.485 ;
        RECT 66.690 1.410 66.970 8.485 ;
        RECT 68.690 1.410 70.335 8.805 ;
        RECT 72.055 1.410 111.095 8.805 ;
        RECT 112.815 8.485 118.675 8.805 ;
        RECT 112.815 1.410 116.720 8.485 ;
        RECT 118.440 1.410 118.675 8.485 ;
        RECT 120.395 16.915 153.995 17.210 ;
        RECT 120.395 1.410 139.380 16.915 ;
        RECT 141.100 15.320 153.995 16.915 ;
        RECT 141.100 12.920 148.225 15.320 ;
        RECT 141.100 1.410 144.730 12.920 ;
        RECT 146.450 1.410 148.225 12.920 ;
        RECT 149.945 1.410 153.995 15.320 ;
        RECT 155.715 1.410 162.460 29.895 ;
        RECT 164.180 1.410 170.915 29.895 ;
        RECT 172.635 16.450 251.410 29.895 ;
        RECT 172.635 1.410 202.640 16.450 ;
        RECT 204.360 1.410 251.410 16.450 ;
        RECT 253.130 25.975 430.450 36.690 ;
        RECT 253.130 18.945 306.935 25.975 ;
        RECT 253.130 17.655 281.025 18.945 ;
        RECT 253.130 1.410 268.560 17.655 ;
        RECT 270.280 15.420 281.025 17.655 ;
        RECT 270.280 1.410 271.785 15.420 ;
        RECT 273.505 13.000 281.025 15.420 ;
        RECT 273.505 1.410 275.520 13.000 ;
        RECT 277.240 1.410 281.025 13.000 ;
        RECT 282.745 1.410 306.935 18.945 ;
        RECT 308.655 8.805 416.560 25.975 ;
        RECT 308.655 8.485 314.490 8.805 ;
        RECT 308.655 1.410 310.275 8.485 ;
        RECT 311.995 1.410 314.490 8.485 ;
        RECT 316.210 1.410 355.245 8.805 ;
        RECT 356.965 1.410 358.610 8.805 ;
        RECT 360.330 8.485 364.850 8.805 ;
        RECT 360.330 1.410 360.600 8.485 ;
        RECT 362.320 1.410 362.850 8.485 ;
        RECT 364.570 1.410 364.850 8.485 ;
        RECT 366.570 1.410 368.215 8.805 ;
        RECT 369.935 1.410 408.975 8.805 ;
        RECT 410.695 8.485 416.560 8.805 ;
        RECT 410.695 1.410 413.175 8.485 ;
        RECT 414.895 1.410 416.560 8.485 ;
        RECT 418.280 1.410 430.450 25.975 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 431.860 484.880 ;
  END
END gf180_ram_512x8_wrapper
END LIBRARY

