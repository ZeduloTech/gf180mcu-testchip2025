VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2900.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 11.080 11.440 20.080 988.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 11.080 11.440 2887.480 20.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 11.080 979.160 2887.480 988.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2878.480 11.440 2887.480 988.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.330 0.440 28.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.330 0.440 108.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.330 0.440 188.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.330 0.440 268.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.330 0.440 348.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.330 0.440 428.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.330 0.440 508.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.330 0.440 588.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.330 0.440 668.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.330 0.440 748.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.330 0.440 828.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.330 0.440 908.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.330 0.440 988.830 79.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.330 578.440 988.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.330 0.440 1068.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.330 0.440 1148.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.330 0.440 1228.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.330 0.440 1308.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.330 0.440 1388.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.330 0.440 1468.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.330 0.440 1548.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.330 0.440 1628.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.330 0.440 1708.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.330 0.440 1788.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.330 0.440 1868.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.330 0.440 1948.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.330 0.440 2028.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.330 0.440 2108.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.330 0.440 2188.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.330 0.440 2268.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.330 0.440 2348.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.330 0.440 2428.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.330 0.440 2508.830 96.330 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.330 184.390 2508.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.330 0.440 2588.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.330 0.440 2668.830 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.330 144.725 2668.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.330 0.440 2748.830 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.330 0.440 2828.830 999.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 56.840 2898.480 59.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 116.840 2635.895 119.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 176.840 2898.480 179.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 236.840 2898.480 239.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 296.840 2898.480 299.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 356.840 2898.480 359.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 416.840 2898.480 419.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 476.840 2898.480 479.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 536.840 2898.480 539.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 596.840 2898.480 599.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 656.840 2898.480 659.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 716.840 2898.480 719.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 776.840 2898.480 779.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 836.840 2898.480 839.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 896.840 2898.480 899.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 956.840 2898.480 959.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 116.840 2898.480 119.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2620.830 0.440 2623.330 999.160 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.080 0.440 9.080 999.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 0.440 2898.480 9.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 990.160 2898.480 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2889.480 0.440 2898.480 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 47.830 0.440 50.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.830 0.440 130.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.830 0.440 210.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 287.830 0.440 290.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 367.830 0.440 370.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 447.830 0.440 450.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 527.830 0.440 530.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 607.830 0.440 610.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 687.830 0.440 690.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 767.830 0.440 770.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 847.830 0.440 850.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 927.830 0.440 930.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1007.830 0.440 1010.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1087.830 0.440 1090.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1167.830 0.440 1170.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1247.830 0.440 1250.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.830 0.440 1330.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1407.830 0.440 1410.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1487.830 0.440 1490.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1567.830 0.440 1570.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1647.830 0.440 1650.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1727.830 0.440 1730.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1807.830 0.440 1810.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1887.830 0.440 1890.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1967.830 0.440 1970.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2047.830 0.440 2050.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2127.830 0.440 2130.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2207.830 0.440 2210.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.830 0.440 2290.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2367.830 0.440 2370.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2447.830 0.440 2450.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2527.830 0.440 2530.330 96.330 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2527.830 184.390 2530.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2607.830 0.440 2610.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2687.830 0.440 2690.330 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2687.830 144.725 2690.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2767.830 0.440 2770.330 999.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2847.830 0.440 2850.330 999.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 86.340 2636.395 88.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 146.340 2635.895 148.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 206.340 2898.480 208.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 266.340 2898.480 268.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 326.340 2898.480 328.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 386.340 2898.480 388.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 446.340 2898.480 448.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 506.340 2898.480 508.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 566.340 2898.480 568.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 626.340 2898.480 628.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 686.340 2898.480 688.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 746.340 2898.480 748.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 806.340 2898.480 808.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 866.340 2898.480 868.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.080 926.340 2898.480 928.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 86.340 2898.480 88.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2707.455 146.340 2898.480 148.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2632.330 0.440 2634.830 999.160 ;
    END
  END VSS
  PIN caravel_io_ie[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 0.000 91.560 1.120 ;
    END
  END caravel_io_ie[0]
  PIN caravel_io_ie[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2240.840 0.000 2241.960 1.120 ;
    END
  END caravel_io_ie[10]
  PIN caravel_io_ie[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2455.880 0.000 2457.000 1.120 ;
    END
  END caravel_io_ie[11]
  PIN caravel_io_ie[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2670.920 0.000 2672.040 1.120 ;
    END
  END caravel_io_ie[12]
  PIN caravel_io_ie[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 305.480 0.000 306.600 1.120 ;
    END
  END caravel_io_ie[1]
  PIN caravel_io_ie[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 520.520 0.000 521.640 1.120 ;
    END
  END caravel_io_ie[2]
  PIN caravel_io_ie[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 735.560 0.000 736.680 1.120 ;
    END
  END caravel_io_ie[3]
  PIN caravel_io_ie[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 950.600 0.000 951.720 1.120 ;
    END
  END caravel_io_ie[4]
  PIN caravel_io_ie[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.640 0.000 1166.760 1.120 ;
    END
  END caravel_io_ie[5]
  PIN caravel_io_ie[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.680 0.000 1381.800 1.120 ;
    END
  END caravel_io_ie[6]
  PIN caravel_io_ie[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1595.720 0.000 1596.840 1.120 ;
    END
  END caravel_io_ie[7]
  PIN caravel_io_ie[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1810.760 0.000 1811.880 1.120 ;
    END
  END caravel_io_ie[8]
  PIN caravel_io_ie[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2025.800 0.000 2026.920 1.120 ;
    END
  END caravel_io_ie[9]
  PIN caravel_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.320 0.000 118.440 1.120 ;
    END
  END caravel_io_in[0]
  PIN caravel_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2267.720 0.000 2268.840 1.120 ;
    END
  END caravel_io_in[10]
  PIN caravel_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2482.760 0.000 2483.880 1.120 ;
    END
  END caravel_io_in[11]
  PIN caravel_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.573000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 2697.800 0.000 2698.920 1.120 ;
    END
  END caravel_io_in[12]
  PIN caravel_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 332.360 0.000 333.480 1.120 ;
    END
  END caravel_io_in[1]
  PIN caravel_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.400 0.000 548.520 1.120 ;
    END
  END caravel_io_in[2]
  PIN caravel_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.440 0.000 763.560 1.120 ;
    END
  END caravel_io_in[3]
  PIN caravel_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.942000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 977.480 0.000 978.600 1.120 ;
    END
  END caravel_io_in[4]
  PIN caravel_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.520 0.000 1193.640 1.120 ;
    END
  END caravel_io_in[5]
  PIN caravel_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1407.560 0.000 1408.680 1.120 ;
    END
  END caravel_io_in[6]
  PIN caravel_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.600 0.000 1623.720 1.120 ;
    END
  END caravel_io_in[7]
  PIN caravel_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.573000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1837.640 0.000 1838.760 1.120 ;
    END
  END caravel_io_in[8]
  PIN caravel_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2052.680 0.000 2053.800 1.120 ;
    END
  END caravel_io_in[9]
  PIN caravel_io_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 0.000 145.320 1.120 ;
    END
  END caravel_io_oe[0]
  PIN caravel_io_oe[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2294.600 0.000 2295.720 1.120 ;
    END
  END caravel_io_oe[10]
  PIN caravel_io_oe[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2509.640 0.000 2510.760 1.120 ;
    END
  END caravel_io_oe[11]
  PIN caravel_io_oe[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2724.680 0.000 2725.800 1.120 ;
    END
  END caravel_io_oe[12]
  PIN caravel_io_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.240 0.000 360.360 1.120 ;
    END
  END caravel_io_oe[1]
  PIN caravel_io_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.280 0.000 575.400 1.120 ;
    END
  END caravel_io_oe[2]
  PIN caravel_io_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 789.320 0.000 790.440 1.120 ;
    END
  END caravel_io_oe[3]
  PIN caravel_io_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.360 0.000 1005.480 1.120 ;
    END
  END caravel_io_oe[4]
  PIN caravel_io_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1219.400 0.000 1220.520 1.120 ;
    END
  END caravel_io_oe[5]
  PIN caravel_io_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.440 0.000 1435.560 1.120 ;
    END
  END caravel_io_oe[6]
  PIN caravel_io_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1649.480 0.000 1650.600 1.120 ;
    END
  END caravel_io_oe[7]
  PIN caravel_io_oe[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1864.520 0.000 1865.640 1.120 ;
    END
  END caravel_io_oe[8]
  PIN caravel_io_oe[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2079.560 0.000 2080.680 1.120 ;
    END
  END caravel_io_oe[9]
  PIN caravel_io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 171.080 0.000 172.200 1.120 ;
    END
  END caravel_io_out[0]
  PIN caravel_io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2321.480 0.000 2322.600 1.120 ;
    END
  END caravel_io_out[10]
  PIN caravel_io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2536.520 0.000 2537.640 1.120 ;
    END
  END caravel_io_out[11]
  PIN caravel_io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2751.560 0.000 2752.680 1.120 ;
    END
  END caravel_io_out[12]
  PIN caravel_io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.120 0.000 387.240 1.120 ;
    END
  END caravel_io_out[1]
  PIN caravel_io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 601.160 0.000 602.280 1.120 ;
    END
  END caravel_io_out[2]
  PIN caravel_io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 816.200 0.000 817.320 1.120 ;
    END
  END caravel_io_out[3]
  PIN caravel_io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.240 0.000 1032.360 1.120 ;
    END
  END caravel_io_out[4]
  PIN caravel_io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1246.280 0.000 1247.400 1.120 ;
    END
  END caravel_io_out[5]
  PIN caravel_io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1461.320 0.000 1462.440 1.120 ;
    END
  END caravel_io_out[6]
  PIN caravel_io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1676.360 0.000 1677.480 1.120 ;
    END
  END caravel_io_out[7]
  PIN caravel_io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1891.400 0.000 1892.520 1.120 ;
    END
  END caravel_io_out[8]
  PIN caravel_io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2106.440 0.000 2107.560 1.120 ;
    END
  END caravel_io_out[9]
  PIN caravel_io_pulldown_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 197.960 0.000 199.080 1.120 ;
    END
  END caravel_io_pulldown_sel[0]
  PIN caravel_io_pulldown_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2348.360 0.000 2349.480 1.120 ;
    END
  END caravel_io_pulldown_sel[10]
  PIN caravel_io_pulldown_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2563.400 0.000 2564.520 1.120 ;
    END
  END caravel_io_pulldown_sel[11]
  PIN caravel_io_pulldown_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2778.440 0.000 2779.560 1.120 ;
    END
  END caravel_io_pulldown_sel[12]
  PIN caravel_io_pulldown_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.000 0.000 414.120 1.120 ;
    END
  END caravel_io_pulldown_sel[1]
  PIN caravel_io_pulldown_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 628.040 0.000 629.160 1.120 ;
    END
  END caravel_io_pulldown_sel[2]
  PIN caravel_io_pulldown_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 843.080 0.000 844.200 1.120 ;
    END
  END caravel_io_pulldown_sel[3]
  PIN caravel_io_pulldown_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.120 0.000 1059.240 1.120 ;
    END
  END caravel_io_pulldown_sel[4]
  PIN caravel_io_pulldown_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.160 0.000 1274.280 1.120 ;
    END
  END caravel_io_pulldown_sel[5]
  PIN caravel_io_pulldown_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1488.200 0.000 1489.320 1.120 ;
    END
  END caravel_io_pulldown_sel[6]
  PIN caravel_io_pulldown_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1703.240 0.000 1704.360 1.120 ;
    END
  END caravel_io_pulldown_sel[7]
  PIN caravel_io_pulldown_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1918.280 0.000 1919.400 1.120 ;
    END
  END caravel_io_pulldown_sel[8]
  PIN caravel_io_pulldown_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2133.320 0.000 2134.440 1.120 ;
    END
  END caravel_io_pulldown_sel[9]
  PIN caravel_io_pullup_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 224.840 0.000 225.960 1.120 ;
    END
  END caravel_io_pullup_sel[0]
  PIN caravel_io_pullup_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2375.240 0.000 2376.360 1.120 ;
    END
  END caravel_io_pullup_sel[10]
  PIN caravel_io_pullup_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2590.280 0.000 2591.400 1.120 ;
    END
  END caravel_io_pullup_sel[11]
  PIN caravel_io_pullup_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2805.320 0.000 2806.440 1.120 ;
    END
  END caravel_io_pullup_sel[12]
  PIN caravel_io_pullup_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 439.880 0.000 441.000 1.120 ;
    END
  END caravel_io_pullup_sel[1]
  PIN caravel_io_pullup_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 654.920 0.000 656.040 1.120 ;
    END
  END caravel_io_pullup_sel[2]
  PIN caravel_io_pullup_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 869.960 0.000 871.080 1.120 ;
    END
  END caravel_io_pullup_sel[3]
  PIN caravel_io_pullup_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1085.000 0.000 1086.120 1.120 ;
    END
  END caravel_io_pullup_sel[4]
  PIN caravel_io_pullup_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.040 0.000 1301.160 1.120 ;
    END
  END caravel_io_pullup_sel[5]
  PIN caravel_io_pullup_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.080 0.000 1516.200 1.120 ;
    END
  END caravel_io_pullup_sel[6]
  PIN caravel_io_pullup_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1730.120 0.000 1731.240 1.120 ;
    END
  END caravel_io_pullup_sel[7]
  PIN caravel_io_pullup_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1945.160 0.000 1946.280 1.120 ;
    END
  END caravel_io_pullup_sel[8]
  PIN caravel_io_pullup_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2160.200 0.000 2161.320 1.120 ;
    END
  END caravel_io_pullup_sel[9]
  PIN caravel_io_schmitt_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 251.720 0.000 252.840 1.120 ;
    END
  END caravel_io_schmitt_sel[0]
  PIN caravel_io_schmitt_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2402.120 0.000 2403.240 1.120 ;
    END
  END caravel_io_schmitt_sel[10]
  PIN caravel_io_schmitt_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2617.160 0.000 2618.280 1.120 ;
    END
  END caravel_io_schmitt_sel[11]
  PIN caravel_io_schmitt_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2832.200 0.000 2833.320 1.120 ;
    END
  END caravel_io_schmitt_sel[12]
  PIN caravel_io_schmitt_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 466.760 0.000 467.880 1.120 ;
    END
  END caravel_io_schmitt_sel[1]
  PIN caravel_io_schmitt_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 681.800 0.000 682.920 1.120 ;
    END
  END caravel_io_schmitt_sel[2]
  PIN caravel_io_schmitt_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 896.840 0.000 897.960 1.120 ;
    END
  END caravel_io_schmitt_sel[3]
  PIN caravel_io_schmitt_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1111.880 0.000 1113.000 1.120 ;
    END
  END caravel_io_schmitt_sel[4]
  PIN caravel_io_schmitt_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1326.920 0.000 1328.040 1.120 ;
    END
  END caravel_io_schmitt_sel[5]
  PIN caravel_io_schmitt_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1541.960 0.000 1543.080 1.120 ;
    END
  END caravel_io_schmitt_sel[6]
  PIN caravel_io_schmitt_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.000 0.000 1758.120 1.120 ;
    END
  END caravel_io_schmitt_sel[7]
  PIN caravel_io_schmitt_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1972.040 0.000 1973.160 1.120 ;
    END
  END caravel_io_schmitt_sel[8]
  PIN caravel_io_schmitt_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2187.080 0.000 2188.200 1.120 ;
    END
  END caravel_io_schmitt_sel[9]
  PIN caravel_io_slew_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 0.000 279.720 1.120 ;
    END
  END caravel_io_slew_sel[0]
  PIN caravel_io_slew_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2429.000 0.000 2430.120 1.120 ;
    END
  END caravel_io_slew_sel[10]
  PIN caravel_io_slew_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2644.040 0.000 2645.160 1.120 ;
    END
  END caravel_io_slew_sel[11]
  PIN caravel_io_slew_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2859.080 0.000 2860.200 1.120 ;
    END
  END caravel_io_slew_sel[12]
  PIN caravel_io_slew_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 493.640 0.000 494.760 1.120 ;
    END
  END caravel_io_slew_sel[1]
  PIN caravel_io_slew_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 708.680 0.000 709.800 1.120 ;
    END
  END caravel_io_slew_sel[2]
  PIN caravel_io_slew_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 923.720 0.000 924.840 1.120 ;
    END
  END caravel_io_slew_sel[3]
  PIN caravel_io_slew_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1138.760 0.000 1139.880 1.120 ;
    END
  END caravel_io_slew_sel[4]
  PIN caravel_io_slew_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1353.800 0.000 1354.920 1.120 ;
    END
  END caravel_io_slew_sel[5]
  PIN caravel_io_slew_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1568.840 0.000 1569.960 1.120 ;
    END
  END caravel_io_slew_sel[6]
  PIN caravel_io_slew_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1783.880 0.000 1785.000 1.120 ;
    END
  END caravel_io_slew_sel[7]
  PIN caravel_io_slew_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1998.920 0.000 2000.040 1.120 ;
    END
  END caravel_io_slew_sel[8]
  PIN caravel_io_slew_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2213.960 0.000 2215.080 1.120 ;
    END
  END caravel_io_slew_sel[9]
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.680 0.000 37.800 1.120 ;
    END
  END clock_core
  PIN flash_clk_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.130000 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 404.600 2900.000 405.720 ;
    END
  END flash_clk_frame
  PIN flash_clk_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 466.760 2900.000 467.880 ;
    END
  END flash_clk_oe
  PIN flash_csb_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 280.280 2900.000 281.400 ;
    END
  END flash_csb_frame
  PIN flash_csb_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 342.440 2900.000 343.560 ;
    END
  END flash_csb_oe
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 528.920 2900.000 530.040 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 591.080 2900.000 592.200 ;
    END
  END flash_io0_do
  PIN flash_io0_ie
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 653.240 2900.000 654.360 ;
    END
  END flash_io0_ie
  PIN flash_io0_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 715.400 2900.000 716.520 ;
    END
  END flash_io0_oe
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 777.560 2900.000 778.680 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 839.720 2900.000 840.840 ;
    END
  END flash_io1_do
  PIN flash_io1_ie
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 901.880 2900.000 903.000 ;
    END
  END flash_io1_ie
  PIN flash_io1_oe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 964.040 2900.000 965.160 ;
    END
  END flash_io1_oe
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 31.640 2900.000 32.760 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 93.800 2900.000 94.920 ;
    END
  END gpio_inenb_core
  PIN gpio_out_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 155.960 2900.000 157.080 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2898.880 218.120 2900.000 219.240 ;
    END
  END gpio_outenb_core
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.560 0.000 64.680 1.120 ;
    END
  END rstb
  PIN user_clock2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2076.200 998.880 2077.320 1000.000 ;
    END
  END user_clock2
  PIN user_gpio_in[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2094.680 998.880 2095.800 1000.000 ;
    END
  END user_gpio_in[0]
  PIN user_gpio_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2649.080 998.880 2650.200 1000.000 ;
    END
  END user_gpio_in[10]
  PIN user_gpio_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2704.520 998.880 2705.640 1000.000 ;
    END
  END user_gpio_in[11]
  PIN user_gpio_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2759.960 998.880 2761.080 1000.000 ;
    END
  END user_gpio_in[12]
  PIN user_gpio_in[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2150.120 998.880 2151.240 1000.000 ;
    END
  END user_gpio_in[1]
  PIN user_gpio_in[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2205.560 998.880 2206.680 1000.000 ;
    END
  END user_gpio_in[2]
  PIN user_gpio_in[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2261.000 998.880 2262.120 1000.000 ;
    END
  END user_gpio_in[3]
  PIN user_gpio_in[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2316.440 998.880 2317.560 1000.000 ;
    END
  END user_gpio_in[4]
  PIN user_gpio_in[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2371.880 998.880 2373.000 1000.000 ;
    END
  END user_gpio_in[5]
  PIN user_gpio_in[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2427.320 998.880 2428.440 1000.000 ;
    END
  END user_gpio_in[6]
  PIN user_gpio_in[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2482.760 998.880 2483.880 1000.000 ;
    END
  END user_gpio_in[7]
  PIN user_gpio_in[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2538.200 998.880 2539.320 1000.000 ;
    END
  END user_gpio_in[8]
  PIN user_gpio_in[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2593.640 998.880 2594.760 1000.000 ;
    END
  END user_gpio_in[9]
  PIN user_gpio_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2113.160 998.880 2114.280 1000.000 ;
    END
  END user_gpio_oeb[0]
  PIN user_gpio_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2667.560 998.880 2668.680 1000.000 ;
    END
  END user_gpio_oeb[10]
  PIN user_gpio_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2723.000 998.880 2724.120 1000.000 ;
    END
  END user_gpio_oeb[11]
  PIN user_gpio_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2778.440 998.880 2779.560 1000.000 ;
    END
  END user_gpio_oeb[12]
  PIN user_gpio_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2168.600 998.880 2169.720 1000.000 ;
    END
  END user_gpio_oeb[1]
  PIN user_gpio_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2224.040 998.880 2225.160 1000.000 ;
    END
  END user_gpio_oeb[2]
  PIN user_gpio_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2279.480 998.880 2280.600 1000.000 ;
    END
  END user_gpio_oeb[3]
  PIN user_gpio_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2334.920 998.880 2336.040 1000.000 ;
    END
  END user_gpio_oeb[4]
  PIN user_gpio_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2390.360 998.880 2391.480 1000.000 ;
    END
  END user_gpio_oeb[5]
  PIN user_gpio_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2445.800 998.880 2446.920 1000.000 ;
    END
  END user_gpio_oeb[6]
  PIN user_gpio_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2501.240 998.880 2502.360 1000.000 ;
    END
  END user_gpio_oeb[7]
  PIN user_gpio_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2556.680 998.880 2557.800 1000.000 ;
    END
  END user_gpio_oeb[8]
  PIN user_gpio_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2612.120 998.880 2613.240 1000.000 ;
    END
  END user_gpio_oeb[9]
  PIN user_gpio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2131.640 998.880 2132.760 1000.000 ;
    END
  END user_gpio_out[0]
  PIN user_gpio_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2686.040 998.880 2687.160 1000.000 ;
    END
  END user_gpio_out[10]
  PIN user_gpio_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2741.480 998.880 2742.600 1000.000 ;
    END
  END user_gpio_out[11]
  PIN user_gpio_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2796.920 998.880 2798.040 1000.000 ;
    END
  END user_gpio_out[12]
  PIN user_gpio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2187.080 998.880 2188.200 1000.000 ;
    END
  END user_gpio_out[1]
  PIN user_gpio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2242.520 998.880 2243.640 1000.000 ;
    END
  END user_gpio_out[2]
  PIN user_gpio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2297.960 998.880 2299.080 1000.000 ;
    END
  END user_gpio_out[3]
  PIN user_gpio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2353.400 998.880 2354.520 1000.000 ;
    END
  END user_gpio_out[4]
  PIN user_gpio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2408.840 998.880 2409.960 1000.000 ;
    END
  END user_gpio_out[5]
  PIN user_gpio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2464.280 998.880 2465.400 1000.000 ;
    END
  END user_gpio_out[6]
  PIN user_gpio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2519.720 998.880 2520.840 1000.000 ;
    END
  END user_gpio_out[7]
  PIN user_gpio_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2575.160 998.880 2576.280 1000.000 ;
    END
  END user_gpio_out[8]
  PIN user_gpio_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2630.600 998.880 2631.720 1000.000 ;
    END
  END user_gpio_out[9]
  PIN user_irq_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2057.720 998.880 2058.840 1000.000 ;
    END
  END user_irq_core
  PIN user_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2020.760 998.880 2021.880 1000.000 ;
    END
  END user_wb_ack_i
  PIN user_wb_adr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 172.760 998.880 173.880 1000.000 ;
    END
  END user_wb_adr_o[0]
  PIN user_wb_adr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 357.560 998.880 358.680 1000.000 ;
    END
  END user_wb_adr_o[10]
  PIN user_wb_adr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 376.040 998.880 377.160 1000.000 ;
    END
  END user_wb_adr_o[11]
  PIN user_wb_adr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 394.520 998.880 395.640 1000.000 ;
    END
  END user_wb_adr_o[12]
  PIN user_wb_adr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.000 998.880 414.120 1000.000 ;
    END
  END user_wb_adr_o[13]
  PIN user_wb_adr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 431.480 998.880 432.600 1000.000 ;
    END
  END user_wb_adr_o[14]
  PIN user_wb_adr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 449.960 998.880 451.080 1000.000 ;
    END
  END user_wb_adr_o[15]
  PIN user_wb_adr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 468.440 998.880 469.560 1000.000 ;
    END
  END user_wb_adr_o[16]
  PIN user_wb_adr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 486.920 998.880 488.040 1000.000 ;
    END
  END user_wb_adr_o[17]
  PIN user_wb_adr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 505.400 998.880 506.520 1000.000 ;
    END
  END user_wb_adr_o[18]
  PIN user_wb_adr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 523.880 998.880 525.000 1000.000 ;
    END
  END user_wb_adr_o[19]
  PIN user_wb_adr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 998.880 192.360 1000.000 ;
    END
  END user_wb_adr_o[1]
  PIN user_wb_adr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 542.360 998.880 543.480 1000.000 ;
    END
  END user_wb_adr_o[20]
  PIN user_wb_adr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 560.840 998.880 561.960 1000.000 ;
    END
  END user_wb_adr_o[21]
  PIN user_wb_adr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 579.320 998.880 580.440 1000.000 ;
    END
  END user_wb_adr_o[22]
  PIN user_wb_adr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 597.800 998.880 598.920 1000.000 ;
    END
  END user_wb_adr_o[23]
  PIN user_wb_adr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 616.280 998.880 617.400 1000.000 ;
    END
  END user_wb_adr_o[24]
  PIN user_wb_adr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 634.760 998.880 635.880 1000.000 ;
    END
  END user_wb_adr_o[25]
  PIN user_wb_adr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 653.240 998.880 654.360 1000.000 ;
    END
  END user_wb_adr_o[26]
  PIN user_wb_adr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 671.720 998.880 672.840 1000.000 ;
    END
  END user_wb_adr_o[27]
  PIN user_wb_adr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 690.200 998.880 691.320 1000.000 ;
    END
  END user_wb_adr_o[28]
  PIN user_wb_adr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 708.680 998.880 709.800 1000.000 ;
    END
  END user_wb_adr_o[29]
  PIN user_wb_adr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 209.720 998.880 210.840 1000.000 ;
    END
  END user_wb_adr_o[2]
  PIN user_wb_adr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 727.160 998.880 728.280 1000.000 ;
    END
  END user_wb_adr_o[30]
  PIN user_wb_adr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 745.640 998.880 746.760 1000.000 ;
    END
  END user_wb_adr_o[31]
  PIN user_wb_adr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 998.880 229.320 1000.000 ;
    END
  END user_wb_adr_o[3]
  PIN user_wb_adr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 246.680 998.880 247.800 1000.000 ;
    END
  END user_wb_adr_o[4]
  PIN user_wb_adr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.160 998.880 266.280 1000.000 ;
    END
  END user_wb_adr_o[5]
  PIN user_wb_adr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 283.640 998.880 284.760 1000.000 ;
    END
  END user_wb_adr_o[6]
  PIN user_wb_adr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 302.120 998.880 303.240 1000.000 ;
    END
  END user_wb_adr_o[7]
  PIN user_wb_adr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 320.600 998.880 321.720 1000.000 ;
    END
  END user_wb_adr_o[8]
  PIN user_wb_adr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 339.080 998.880 340.200 1000.000 ;
    END
  END user_wb_adr_o[9]
  PIN user_wb_clk_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.130000 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.240 998.880 2040.360 1000.000 ;
    END
  END user_wb_clk_o
  PIN user_wb_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1965.320 998.880 1966.440 1000.000 ;
    END
  END user_wb_cyc_o
  PIN user_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1355.480 998.880 1356.600 1000.000 ;
    END
  END user_wb_dat_i[0]
  PIN user_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1540.280 998.880 1541.400 1000.000 ;
    END
  END user_wb_dat_i[10]
  PIN user_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1558.760 998.880 1559.880 1000.000 ;
    END
  END user_wb_dat_i[11]
  PIN user_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1577.240 998.880 1578.360 1000.000 ;
    END
  END user_wb_dat_i[12]
  PIN user_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1595.720 998.880 1596.840 1000.000 ;
    END
  END user_wb_dat_i[13]
  PIN user_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1614.200 998.880 1615.320 1000.000 ;
    END
  END user_wb_dat_i[14]
  PIN user_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1632.680 998.880 1633.800 1000.000 ;
    END
  END user_wb_dat_i[15]
  PIN user_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1651.160 998.880 1652.280 1000.000 ;
    END
  END user_wb_dat_i[16]
  PIN user_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1669.640 998.880 1670.760 1000.000 ;
    END
  END user_wb_dat_i[17]
  PIN user_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1688.120 998.880 1689.240 1000.000 ;
    END
  END user_wb_dat_i[18]
  PIN user_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1706.600 998.880 1707.720 1000.000 ;
    END
  END user_wb_dat_i[19]
  PIN user_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1373.960 998.880 1375.080 1000.000 ;
    END
  END user_wb_dat_i[1]
  PIN user_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1725.080 998.880 1726.200 1000.000 ;
    END
  END user_wb_dat_i[20]
  PIN user_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1743.560 998.880 1744.680 1000.000 ;
    END
  END user_wb_dat_i[21]
  PIN user_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1762.040 998.880 1763.160 1000.000 ;
    END
  END user_wb_dat_i[22]
  PIN user_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1780.520 998.880 1781.640 1000.000 ;
    END
  END user_wb_dat_i[23]
  PIN user_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1799.000 998.880 1800.120 1000.000 ;
    END
  END user_wb_dat_i[24]
  PIN user_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1817.480 998.880 1818.600 1000.000 ;
    END
  END user_wb_dat_i[25]
  PIN user_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1835.960 998.880 1837.080 1000.000 ;
    END
  END user_wb_dat_i[26]
  PIN user_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1854.440 998.880 1855.560 1000.000 ;
    END
  END user_wb_dat_i[27]
  PIN user_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1872.920 998.880 1874.040 1000.000 ;
    END
  END user_wb_dat_i[28]
  PIN user_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1891.400 998.880 1892.520 1000.000 ;
    END
  END user_wb_dat_i[29]
  PIN user_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1392.440 998.880 1393.560 1000.000 ;
    END
  END user_wb_dat_i[2]
  PIN user_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1909.880 998.880 1911.000 1000.000 ;
    END
  END user_wb_dat_i[30]
  PIN user_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1928.360 998.880 1929.480 1000.000 ;
    END
  END user_wb_dat_i[31]
  PIN user_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1410.920 998.880 1412.040 1000.000 ;
    END
  END user_wb_dat_i[3]
  PIN user_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1429.400 998.880 1430.520 1000.000 ;
    END
  END user_wb_dat_i[4]
  PIN user_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1447.880 998.880 1449.000 1000.000 ;
    END
  END user_wb_dat_i[5]
  PIN user_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1466.360 998.880 1467.480 1000.000 ;
    END
  END user_wb_dat_i[6]
  PIN user_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1484.840 998.880 1485.960 1000.000 ;
    END
  END user_wb_dat_i[7]
  PIN user_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1503.320 998.880 1504.440 1000.000 ;
    END
  END user_wb_dat_i[8]
  PIN user_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1521.800 998.880 1522.920 1000.000 ;
    END
  END user_wb_dat_i[9]
  PIN user_wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 764.120 998.880 765.240 1000.000 ;
    END
  END user_wb_dat_o[0]
  PIN user_wb_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 948.920 998.880 950.040 1000.000 ;
    END
  END user_wb_dat_o[10]
  PIN user_wb_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 967.400 998.880 968.520 1000.000 ;
    END
  END user_wb_dat_o[11]
  PIN user_wb_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 985.880 998.880 987.000 1000.000 ;
    END
  END user_wb_dat_o[12]
  PIN user_wb_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.360 998.880 1005.480 1000.000 ;
    END
  END user_wb_dat_o[13]
  PIN user_wb_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1022.840 998.880 1023.960 1000.000 ;
    END
  END user_wb_dat_o[14]
  PIN user_wb_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1041.320 998.880 1042.440 1000.000 ;
    END
  END user_wb_dat_o[15]
  PIN user_wb_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1059.800 998.880 1060.920 1000.000 ;
    END
  END user_wb_dat_o[16]
  PIN user_wb_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1078.280 998.880 1079.400 1000.000 ;
    END
  END user_wb_dat_o[17]
  PIN user_wb_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1096.760 998.880 1097.880 1000.000 ;
    END
  END user_wb_dat_o[18]
  PIN user_wb_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1115.240 998.880 1116.360 1000.000 ;
    END
  END user_wb_dat_o[19]
  PIN user_wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 782.600 998.880 783.720 1000.000 ;
    END
  END user_wb_dat_o[1]
  PIN user_wb_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1133.720 998.880 1134.840 1000.000 ;
    END
  END user_wb_dat_o[20]
  PIN user_wb_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.200 998.880 1153.320 1000.000 ;
    END
  END user_wb_dat_o[21]
  PIN user_wb_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1170.680 998.880 1171.800 1000.000 ;
    END
  END user_wb_dat_o[22]
  PIN user_wb_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1189.160 998.880 1190.280 1000.000 ;
    END
  END user_wb_dat_o[23]
  PIN user_wb_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1207.640 998.880 1208.760 1000.000 ;
    END
  END user_wb_dat_o[24]
  PIN user_wb_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1226.120 998.880 1227.240 1000.000 ;
    END
  END user_wb_dat_o[25]
  PIN user_wb_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1244.600 998.880 1245.720 1000.000 ;
    END
  END user_wb_dat_o[26]
  PIN user_wb_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1263.080 998.880 1264.200 1000.000 ;
    END
  END user_wb_dat_o[27]
  PIN user_wb_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1281.560 998.880 1282.680 1000.000 ;
    END
  END user_wb_dat_o[28]
  PIN user_wb_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.040 998.880 1301.160 1000.000 ;
    END
  END user_wb_dat_o[29]
  PIN user_wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 801.080 998.880 802.200 1000.000 ;
    END
  END user_wb_dat_o[2]
  PIN user_wb_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1318.520 998.880 1319.640 1000.000 ;
    END
  END user_wb_dat_o[30]
  PIN user_wb_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1337.000 998.880 1338.120 1000.000 ;
    END
  END user_wb_dat_o[31]
  PIN user_wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 819.560 998.880 820.680 1000.000 ;
    END
  END user_wb_dat_o[3]
  PIN user_wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 838.040 998.880 839.160 1000.000 ;
    END
  END user_wb_dat_o[4]
  PIN user_wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 856.520 998.880 857.640 1000.000 ;
    END
  END user_wb_dat_o[5]
  PIN user_wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 875.000 998.880 876.120 1000.000 ;
    END
  END user_wb_dat_o[6]
  PIN user_wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 893.480 998.880 894.600 1000.000 ;
    END
  END user_wb_dat_o[7]
  PIN user_wb_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 911.960 998.880 913.080 1000.000 ;
    END
  END user_wb_dat_o[8]
  PIN user_wb_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 930.440 998.880 931.560 1000.000 ;
    END
  END user_wb_dat_o[9]
  PIN user_wb_rst_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1946.840 998.880 1947.960 1000.000 ;
    END
  END user_wb_rst_o
  PIN user_wb_sel_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 998.880 99.960 1000.000 ;
    END
  END user_wb_sel_o[0]
  PIN user_wb_sel_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 117.320 998.880 118.440 1000.000 ;
    END
  END user_wb_sel_o[1]
  PIN user_wb_sel_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 135.800 998.880 136.920 1000.000 ;
    END
  END user_wb_sel_o[2]
  PIN user_wb_sel_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 998.880 155.400 1000.000 ;
    END
  END user_wb_sel_o[3]
  PIN user_wb_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1983.800 998.880 1984.920 1000.000 ;
    END
  END user_wb_stb_o
  PIN user_wb_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2002.280 998.880 2003.400 1000.000 ;
    END
  END user_wb_we_o
  OBS
      LAYER Nwell ;
        RECT 23.650 27.010 2874.910 972.590 ;
      LAYER Metal1 ;
        RECT 24.080 27.140 2874.480 972.460 ;
      LAYER Metal2 ;
        RECT 25.340 998.580 98.540 999.460 ;
        RECT 100.260 998.580 117.020 999.460 ;
        RECT 118.740 998.580 135.500 999.460 ;
        RECT 137.220 998.580 153.980 999.460 ;
        RECT 155.700 998.580 172.460 999.460 ;
        RECT 174.180 998.580 190.940 999.460 ;
        RECT 192.660 998.580 209.420 999.460 ;
        RECT 211.140 998.580 227.900 999.460 ;
        RECT 229.620 998.580 246.380 999.460 ;
        RECT 248.100 998.580 264.860 999.460 ;
        RECT 266.580 998.580 283.340 999.460 ;
        RECT 285.060 998.580 301.820 999.460 ;
        RECT 303.540 998.580 320.300 999.460 ;
        RECT 322.020 998.580 338.780 999.460 ;
        RECT 340.500 998.580 357.260 999.460 ;
        RECT 358.980 998.580 375.740 999.460 ;
        RECT 377.460 998.580 394.220 999.460 ;
        RECT 395.940 998.580 412.700 999.460 ;
        RECT 414.420 998.580 431.180 999.460 ;
        RECT 432.900 998.580 449.660 999.460 ;
        RECT 451.380 998.580 468.140 999.460 ;
        RECT 469.860 998.580 486.620 999.460 ;
        RECT 488.340 998.580 505.100 999.460 ;
        RECT 506.820 998.580 523.580 999.460 ;
        RECT 525.300 998.580 542.060 999.460 ;
        RECT 543.780 998.580 560.540 999.460 ;
        RECT 562.260 998.580 579.020 999.460 ;
        RECT 580.740 998.580 597.500 999.460 ;
        RECT 599.220 998.580 615.980 999.460 ;
        RECT 617.700 998.580 634.460 999.460 ;
        RECT 636.180 998.580 652.940 999.460 ;
        RECT 654.660 998.580 671.420 999.460 ;
        RECT 673.140 998.580 689.900 999.460 ;
        RECT 691.620 998.580 708.380 999.460 ;
        RECT 710.100 998.580 726.860 999.460 ;
        RECT 728.580 998.580 745.340 999.460 ;
        RECT 747.060 998.580 763.820 999.460 ;
        RECT 765.540 998.580 782.300 999.460 ;
        RECT 784.020 998.580 800.780 999.460 ;
        RECT 802.500 998.580 819.260 999.460 ;
        RECT 820.980 998.580 837.740 999.460 ;
        RECT 839.460 998.580 856.220 999.460 ;
        RECT 857.940 998.580 874.700 999.460 ;
        RECT 876.420 998.580 893.180 999.460 ;
        RECT 894.900 998.580 911.660 999.460 ;
        RECT 913.380 998.580 930.140 999.460 ;
        RECT 931.860 998.580 948.620 999.460 ;
        RECT 950.340 998.580 967.100 999.460 ;
        RECT 968.820 998.580 985.580 999.460 ;
        RECT 987.300 998.580 1004.060 999.460 ;
        RECT 1005.780 998.580 1022.540 999.460 ;
        RECT 1024.260 998.580 1041.020 999.460 ;
        RECT 1042.740 998.580 1059.500 999.460 ;
        RECT 1061.220 998.580 1077.980 999.460 ;
        RECT 1079.700 998.580 1096.460 999.460 ;
        RECT 1098.180 998.580 1114.940 999.460 ;
        RECT 1116.660 998.580 1133.420 999.460 ;
        RECT 1135.140 998.580 1151.900 999.460 ;
        RECT 1153.620 998.580 1170.380 999.460 ;
        RECT 1172.100 998.580 1188.860 999.460 ;
        RECT 1190.580 998.580 1207.340 999.460 ;
        RECT 1209.060 998.580 1225.820 999.460 ;
        RECT 1227.540 998.580 1244.300 999.460 ;
        RECT 1246.020 998.580 1262.780 999.460 ;
        RECT 1264.500 998.580 1281.260 999.460 ;
        RECT 1282.980 998.580 1299.740 999.460 ;
        RECT 1301.460 998.580 1318.220 999.460 ;
        RECT 1319.940 998.580 1336.700 999.460 ;
        RECT 1338.420 998.580 1355.180 999.460 ;
        RECT 1356.900 998.580 1373.660 999.460 ;
        RECT 1375.380 998.580 1392.140 999.460 ;
        RECT 1393.860 998.580 1410.620 999.460 ;
        RECT 1412.340 998.580 1429.100 999.460 ;
        RECT 1430.820 998.580 1447.580 999.460 ;
        RECT 1449.300 998.580 1466.060 999.460 ;
        RECT 1467.780 998.580 1484.540 999.460 ;
        RECT 1486.260 998.580 1503.020 999.460 ;
        RECT 1504.740 998.580 1521.500 999.460 ;
        RECT 1523.220 998.580 1539.980 999.460 ;
        RECT 1541.700 998.580 1558.460 999.460 ;
        RECT 1560.180 998.580 1576.940 999.460 ;
        RECT 1578.660 998.580 1595.420 999.460 ;
        RECT 1597.140 998.580 1613.900 999.460 ;
        RECT 1615.620 998.580 1632.380 999.460 ;
        RECT 1634.100 998.580 1650.860 999.460 ;
        RECT 1652.580 998.580 1669.340 999.460 ;
        RECT 1671.060 998.580 1687.820 999.460 ;
        RECT 1689.540 998.580 1706.300 999.460 ;
        RECT 1708.020 998.580 1724.780 999.460 ;
        RECT 1726.500 998.580 1743.260 999.460 ;
        RECT 1744.980 998.580 1761.740 999.460 ;
        RECT 1763.460 998.580 1780.220 999.460 ;
        RECT 1781.940 998.580 1798.700 999.460 ;
        RECT 1800.420 998.580 1817.180 999.460 ;
        RECT 1818.900 998.580 1835.660 999.460 ;
        RECT 1837.380 998.580 1854.140 999.460 ;
        RECT 1855.860 998.580 1872.620 999.460 ;
        RECT 1874.340 998.580 1891.100 999.460 ;
        RECT 1892.820 998.580 1909.580 999.460 ;
        RECT 1911.300 998.580 1928.060 999.460 ;
        RECT 1929.780 998.580 1946.540 999.460 ;
        RECT 1948.260 998.580 1965.020 999.460 ;
        RECT 1966.740 998.580 1983.500 999.460 ;
        RECT 1985.220 998.580 2001.980 999.460 ;
        RECT 2003.700 998.580 2020.460 999.460 ;
        RECT 2022.180 998.580 2038.940 999.460 ;
        RECT 2040.660 998.580 2057.420 999.460 ;
        RECT 2059.140 998.580 2075.900 999.460 ;
        RECT 2077.620 998.580 2094.380 999.460 ;
        RECT 2096.100 998.580 2112.860 999.460 ;
        RECT 2114.580 998.580 2131.340 999.460 ;
        RECT 2133.060 998.580 2149.820 999.460 ;
        RECT 2151.540 998.580 2168.300 999.460 ;
        RECT 2170.020 998.580 2186.780 999.460 ;
        RECT 2188.500 998.580 2205.260 999.460 ;
        RECT 2206.980 998.580 2223.740 999.460 ;
        RECT 2225.460 998.580 2242.220 999.460 ;
        RECT 2243.940 998.580 2260.700 999.460 ;
        RECT 2262.420 998.580 2279.180 999.460 ;
        RECT 2280.900 998.580 2297.660 999.460 ;
        RECT 2299.380 998.580 2316.140 999.460 ;
        RECT 2317.860 998.580 2334.620 999.460 ;
        RECT 2336.340 998.580 2353.100 999.460 ;
        RECT 2354.820 998.580 2371.580 999.460 ;
        RECT 2373.300 998.580 2390.060 999.460 ;
        RECT 2391.780 998.580 2408.540 999.460 ;
        RECT 2410.260 998.580 2427.020 999.460 ;
        RECT 2428.740 998.580 2445.500 999.460 ;
        RECT 2447.220 998.580 2463.980 999.460 ;
        RECT 2465.700 998.580 2482.460 999.460 ;
        RECT 2484.180 998.580 2500.940 999.460 ;
        RECT 2502.660 998.580 2519.420 999.460 ;
        RECT 2521.140 998.580 2537.900 999.460 ;
        RECT 2539.620 998.580 2556.380 999.460 ;
        RECT 2558.100 998.580 2574.860 999.460 ;
        RECT 2576.580 998.580 2593.340 999.460 ;
        RECT 2595.060 998.580 2611.820 999.460 ;
        RECT 2613.540 998.580 2630.300 999.460 ;
        RECT 2632.020 998.580 2648.780 999.460 ;
        RECT 2650.500 998.580 2667.260 999.460 ;
        RECT 2668.980 998.580 2685.740 999.460 ;
        RECT 2687.460 998.580 2704.220 999.460 ;
        RECT 2705.940 998.580 2722.700 999.460 ;
        RECT 2724.420 998.580 2741.180 999.460 ;
        RECT 2742.900 998.580 2759.660 999.460 ;
        RECT 2761.380 998.580 2778.140 999.460 ;
        RECT 2779.860 998.580 2796.620 999.460 ;
        RECT 2798.340 998.580 2872.660 999.460 ;
        RECT 25.340 1.420 2872.660 998.580 ;
        RECT 25.340 0.650 36.380 1.420 ;
        RECT 38.100 0.650 63.260 1.420 ;
        RECT 64.980 0.650 90.140 1.420 ;
        RECT 91.860 0.650 117.020 1.420 ;
        RECT 118.740 0.650 143.900 1.420 ;
        RECT 145.620 0.650 170.780 1.420 ;
        RECT 172.500 0.650 197.660 1.420 ;
        RECT 199.380 0.650 224.540 1.420 ;
        RECT 226.260 0.650 251.420 1.420 ;
        RECT 253.140 0.650 278.300 1.420 ;
        RECT 280.020 0.650 305.180 1.420 ;
        RECT 306.900 0.650 332.060 1.420 ;
        RECT 333.780 0.650 358.940 1.420 ;
        RECT 360.660 0.650 385.820 1.420 ;
        RECT 387.540 0.650 412.700 1.420 ;
        RECT 414.420 0.650 439.580 1.420 ;
        RECT 441.300 0.650 466.460 1.420 ;
        RECT 468.180 0.650 493.340 1.420 ;
        RECT 495.060 0.650 520.220 1.420 ;
        RECT 521.940 0.650 547.100 1.420 ;
        RECT 548.820 0.650 573.980 1.420 ;
        RECT 575.700 0.650 600.860 1.420 ;
        RECT 602.580 0.650 627.740 1.420 ;
        RECT 629.460 0.650 654.620 1.420 ;
        RECT 656.340 0.650 681.500 1.420 ;
        RECT 683.220 0.650 708.380 1.420 ;
        RECT 710.100 0.650 735.260 1.420 ;
        RECT 736.980 0.650 762.140 1.420 ;
        RECT 763.860 0.650 789.020 1.420 ;
        RECT 790.740 0.650 815.900 1.420 ;
        RECT 817.620 0.650 842.780 1.420 ;
        RECT 844.500 0.650 869.660 1.420 ;
        RECT 871.380 0.650 896.540 1.420 ;
        RECT 898.260 0.650 923.420 1.420 ;
        RECT 925.140 0.650 950.300 1.420 ;
        RECT 952.020 0.650 977.180 1.420 ;
        RECT 978.900 0.650 1004.060 1.420 ;
        RECT 1005.780 0.650 1030.940 1.420 ;
        RECT 1032.660 0.650 1057.820 1.420 ;
        RECT 1059.540 0.650 1084.700 1.420 ;
        RECT 1086.420 0.650 1111.580 1.420 ;
        RECT 1113.300 0.650 1138.460 1.420 ;
        RECT 1140.180 0.650 1165.340 1.420 ;
        RECT 1167.060 0.650 1192.220 1.420 ;
        RECT 1193.940 0.650 1219.100 1.420 ;
        RECT 1220.820 0.650 1245.980 1.420 ;
        RECT 1247.700 0.650 1272.860 1.420 ;
        RECT 1274.580 0.650 1299.740 1.420 ;
        RECT 1301.460 0.650 1326.620 1.420 ;
        RECT 1328.340 0.650 1353.500 1.420 ;
        RECT 1355.220 0.650 1380.380 1.420 ;
        RECT 1382.100 0.650 1407.260 1.420 ;
        RECT 1408.980 0.650 1434.140 1.420 ;
        RECT 1435.860 0.650 1461.020 1.420 ;
        RECT 1462.740 0.650 1487.900 1.420 ;
        RECT 1489.620 0.650 1514.780 1.420 ;
        RECT 1516.500 0.650 1541.660 1.420 ;
        RECT 1543.380 0.650 1568.540 1.420 ;
        RECT 1570.260 0.650 1595.420 1.420 ;
        RECT 1597.140 0.650 1622.300 1.420 ;
        RECT 1624.020 0.650 1649.180 1.420 ;
        RECT 1650.900 0.650 1676.060 1.420 ;
        RECT 1677.780 0.650 1702.940 1.420 ;
        RECT 1704.660 0.650 1729.820 1.420 ;
        RECT 1731.540 0.650 1756.700 1.420 ;
        RECT 1758.420 0.650 1783.580 1.420 ;
        RECT 1785.300 0.650 1810.460 1.420 ;
        RECT 1812.180 0.650 1837.340 1.420 ;
        RECT 1839.060 0.650 1864.220 1.420 ;
        RECT 1865.940 0.650 1891.100 1.420 ;
        RECT 1892.820 0.650 1917.980 1.420 ;
        RECT 1919.700 0.650 1944.860 1.420 ;
        RECT 1946.580 0.650 1971.740 1.420 ;
        RECT 1973.460 0.650 1998.620 1.420 ;
        RECT 2000.340 0.650 2025.500 1.420 ;
        RECT 2027.220 0.650 2052.380 1.420 ;
        RECT 2054.100 0.650 2079.260 1.420 ;
        RECT 2080.980 0.650 2106.140 1.420 ;
        RECT 2107.860 0.650 2133.020 1.420 ;
        RECT 2134.740 0.650 2159.900 1.420 ;
        RECT 2161.620 0.650 2186.780 1.420 ;
        RECT 2188.500 0.650 2213.660 1.420 ;
        RECT 2215.380 0.650 2240.540 1.420 ;
        RECT 2242.260 0.650 2267.420 1.420 ;
        RECT 2269.140 0.650 2294.300 1.420 ;
        RECT 2296.020 0.650 2321.180 1.420 ;
        RECT 2322.900 0.650 2348.060 1.420 ;
        RECT 2349.780 0.650 2374.940 1.420 ;
        RECT 2376.660 0.650 2401.820 1.420 ;
        RECT 2403.540 0.650 2428.700 1.420 ;
        RECT 2430.420 0.650 2455.580 1.420 ;
        RECT 2457.300 0.650 2482.460 1.420 ;
        RECT 2484.180 0.650 2509.340 1.420 ;
        RECT 2511.060 0.650 2536.220 1.420 ;
        RECT 2537.940 0.650 2563.100 1.420 ;
        RECT 2564.820 0.650 2589.980 1.420 ;
        RECT 2591.700 0.650 2616.860 1.420 ;
        RECT 2618.580 0.650 2643.740 1.420 ;
        RECT 2645.460 0.650 2670.620 1.420 ;
        RECT 2672.340 0.650 2697.500 1.420 ;
        RECT 2699.220 0.650 2724.380 1.420 ;
        RECT 2726.100 0.650 2751.260 1.420 ;
        RECT 2752.980 0.650 2778.140 1.420 ;
        RECT 2779.860 0.650 2805.020 1.420 ;
        RECT 2806.740 0.650 2831.900 1.420 ;
        RECT 2833.620 0.650 2858.780 1.420 ;
        RECT 2860.500 0.650 2872.660 1.420 ;
      LAYER Metal3 ;
        RECT 25.290 965.460 2899.540 997.220 ;
        RECT 25.290 963.740 2898.580 965.460 ;
        RECT 25.290 903.300 2899.540 963.740 ;
        RECT 25.290 901.580 2898.580 903.300 ;
        RECT 25.290 841.140 2899.540 901.580 ;
        RECT 25.290 839.420 2898.580 841.140 ;
        RECT 25.290 778.980 2899.540 839.420 ;
        RECT 25.290 777.260 2898.580 778.980 ;
        RECT 25.290 716.820 2899.540 777.260 ;
        RECT 25.290 715.100 2898.580 716.820 ;
        RECT 25.290 654.660 2899.540 715.100 ;
        RECT 25.290 652.940 2898.580 654.660 ;
        RECT 25.290 592.500 2899.540 652.940 ;
        RECT 25.290 590.780 2898.580 592.500 ;
        RECT 25.290 530.340 2899.540 590.780 ;
        RECT 25.290 528.620 2898.580 530.340 ;
        RECT 25.290 468.180 2899.540 528.620 ;
        RECT 25.290 466.460 2898.580 468.180 ;
        RECT 25.290 406.020 2899.540 466.460 ;
        RECT 25.290 404.300 2898.580 406.020 ;
        RECT 25.290 343.860 2899.540 404.300 ;
        RECT 25.290 342.140 2898.580 343.860 ;
        RECT 25.290 281.700 2899.540 342.140 ;
        RECT 25.290 279.980 2898.580 281.700 ;
        RECT 25.290 219.540 2899.540 279.980 ;
        RECT 25.290 217.820 2898.580 219.540 ;
        RECT 25.290 157.380 2899.540 217.820 ;
        RECT 25.290 155.660 2898.580 157.380 ;
        RECT 25.290 95.220 2899.540 155.660 ;
        RECT 25.290 93.500 2898.580 95.220 ;
        RECT 25.290 33.060 2899.540 93.500 ;
        RECT 25.290 31.340 2898.580 33.060 ;
        RECT 25.290 0.700 2899.540 31.340 ;
      LAYER Metal4 ;
        RECT 41.580 26.970 47.530 996.150 ;
        RECT 50.630 26.970 106.030 996.150 ;
        RECT 109.130 26.970 127.530 996.150 ;
        RECT 130.630 26.970 186.030 996.150 ;
        RECT 189.130 26.970 207.530 996.150 ;
        RECT 210.630 26.970 266.030 996.150 ;
        RECT 269.130 26.970 287.530 996.150 ;
        RECT 290.630 26.970 346.030 996.150 ;
        RECT 349.130 26.970 367.530 996.150 ;
        RECT 370.630 26.970 426.030 996.150 ;
        RECT 429.130 26.970 447.530 996.150 ;
        RECT 450.630 26.970 506.030 996.150 ;
        RECT 509.130 26.970 527.530 996.150 ;
        RECT 530.630 26.970 586.030 996.150 ;
        RECT 589.130 26.970 607.530 996.150 ;
        RECT 610.630 26.970 666.030 996.150 ;
        RECT 669.130 26.970 687.530 996.150 ;
        RECT 690.630 26.970 746.030 996.150 ;
        RECT 749.130 26.970 767.530 996.150 ;
        RECT 770.630 26.970 826.030 996.150 ;
        RECT 829.130 26.970 847.530 996.150 ;
        RECT 850.630 26.970 906.030 996.150 ;
        RECT 909.130 26.970 927.530 996.150 ;
        RECT 930.630 578.140 986.030 996.150 ;
        RECT 989.130 578.140 1007.530 996.150 ;
        RECT 930.630 79.460 1007.530 578.140 ;
        RECT 930.630 26.970 986.030 79.460 ;
        RECT 989.130 26.970 1007.530 79.460 ;
        RECT 1010.630 26.970 1066.030 996.150 ;
        RECT 1069.130 26.970 1087.530 996.150 ;
        RECT 1090.630 26.970 1146.030 996.150 ;
        RECT 1149.130 26.970 1167.530 996.150 ;
        RECT 1170.630 26.970 1226.030 996.150 ;
        RECT 1229.130 26.970 1247.530 996.150 ;
        RECT 1250.630 26.970 1306.030 996.150 ;
        RECT 1309.130 26.970 1327.530 996.150 ;
        RECT 1330.630 26.970 1386.030 996.150 ;
        RECT 1389.130 26.970 1407.530 996.150 ;
        RECT 1410.630 26.970 1466.030 996.150 ;
        RECT 1469.130 26.970 1487.530 996.150 ;
        RECT 1490.630 26.970 1546.030 996.150 ;
        RECT 1549.130 26.970 1567.530 996.150 ;
        RECT 1570.630 26.970 1626.030 996.150 ;
        RECT 1629.130 26.970 1647.530 996.150 ;
        RECT 1650.630 26.970 1706.030 996.150 ;
        RECT 1709.130 26.970 1727.530 996.150 ;
        RECT 1730.630 26.970 1786.030 996.150 ;
        RECT 1789.130 26.970 1807.530 996.150 ;
        RECT 1810.630 26.970 1866.030 996.150 ;
        RECT 1869.130 26.970 1887.530 996.150 ;
        RECT 1890.630 26.970 1946.030 996.150 ;
        RECT 1949.130 26.970 1967.530 996.150 ;
        RECT 1970.630 26.970 2026.030 996.150 ;
        RECT 2029.130 26.970 2047.530 996.150 ;
        RECT 2050.630 26.970 2106.030 996.150 ;
        RECT 2109.130 26.970 2127.530 996.150 ;
        RECT 2130.630 26.970 2186.030 996.150 ;
        RECT 2189.130 26.970 2207.530 996.150 ;
        RECT 2210.630 26.970 2266.030 996.150 ;
        RECT 2269.130 26.970 2287.530 996.150 ;
        RECT 2290.630 26.970 2346.030 996.150 ;
        RECT 2349.130 26.970 2367.530 996.150 ;
        RECT 2370.630 26.970 2426.030 996.150 ;
        RECT 2429.130 26.970 2447.530 996.150 ;
        RECT 2450.630 184.090 2506.030 996.150 ;
        RECT 2509.130 184.090 2527.530 996.150 ;
        RECT 2530.630 184.090 2586.030 996.150 ;
        RECT 2450.630 96.630 2586.030 184.090 ;
        RECT 2450.630 26.970 2506.030 96.630 ;
        RECT 2509.130 26.970 2527.530 96.630 ;
        RECT 2530.630 26.970 2586.030 96.630 ;
        RECT 2589.130 26.970 2607.530 996.150 ;
        RECT 2610.630 26.970 2620.530 996.150 ;
        RECT 2623.630 26.970 2632.030 996.150 ;
        RECT 2635.130 144.425 2666.030 996.150 ;
        RECT 2669.130 144.425 2687.530 996.150 ;
        RECT 2690.630 144.425 2746.030 996.150 ;
        RECT 2635.130 87.030 2746.030 144.425 ;
        RECT 2635.130 26.970 2666.030 87.030 ;
        RECT 2669.130 26.970 2687.530 87.030 ;
        RECT 2690.630 26.970 2746.030 87.030 ;
        RECT 2749.130 26.970 2767.530 996.150 ;
        RECT 2770.630 26.970 2826.030 996.150 ;
        RECT 2829.130 26.970 2830.100 996.150 ;
      LAYER Metal5 ;
        RECT 154.060 959.940 2792.660 975.370 ;
        RECT 154.060 929.440 2792.660 956.240 ;
        RECT 154.060 899.940 2792.660 925.740 ;
        RECT 154.060 869.440 2792.660 896.240 ;
        RECT 154.060 839.940 2792.660 865.740 ;
        RECT 154.060 809.440 2792.660 836.240 ;
        RECT 154.060 779.940 2792.660 805.740 ;
        RECT 154.060 749.440 2792.660 776.240 ;
        RECT 154.060 719.940 2792.660 745.740 ;
        RECT 154.060 689.440 2792.660 716.240 ;
        RECT 154.060 659.940 2792.660 685.740 ;
        RECT 154.060 629.440 2792.660 656.240 ;
        RECT 154.060 599.940 2792.660 625.740 ;
        RECT 154.060 569.440 2792.660 596.240 ;
        RECT 154.060 539.940 2792.660 565.740 ;
        RECT 154.060 509.440 2792.660 536.240 ;
        RECT 154.060 479.940 2792.660 505.740 ;
        RECT 154.060 449.440 2792.660 476.240 ;
        RECT 154.060 419.940 2792.660 445.740 ;
        RECT 154.060 389.440 2792.660 416.240 ;
        RECT 154.060 359.940 2792.660 385.740 ;
        RECT 154.060 329.440 2792.660 356.240 ;
        RECT 154.060 299.940 2792.660 325.740 ;
        RECT 154.060 269.440 2792.660 296.240 ;
        RECT 154.060 239.940 2792.660 265.740 ;
        RECT 154.060 209.440 2792.660 236.240 ;
        RECT 154.060 179.940 2792.660 205.740 ;
        RECT 154.060 149.440 2792.660 176.240 ;
        RECT 2636.495 145.740 2706.855 149.440 ;
        RECT 154.060 119.940 2792.660 145.740 ;
        RECT 2636.495 116.240 2706.855 119.940 ;
        RECT 154.060 89.440 2792.660 116.240 ;
        RECT 2636.995 85.740 2706.855 89.440 ;
        RECT 154.060 59.940 2792.660 85.740 ;
        RECT 154.060 28.130 2792.660 56.240 ;
  END
END caravel_core
END LIBRARY

