module efuse_wb_mem_1024x32 (wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rst_i,
    wb_stb_i,
    wb_we_i,
    write_enable_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rst_i;
 input wb_stb_i;
 input wb_we_i;
 input write_enable_i;
 input [9:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire \bit_sel[0] ;
 wire \bit_sel[10] ;
 wire \bit_sel[11] ;
 wire \bit_sel[12] ;
 wire \bit_sel[13] ;
 wire \bit_sel[14] ;
 wire \bit_sel[15] ;
 wire \bit_sel[16] ;
 wire \bit_sel[17] ;
 wire \bit_sel[18] ;
 wire \bit_sel[19] ;
 wire \bit_sel[1] ;
 wire \bit_sel[20] ;
 wire \bit_sel[21] ;
 wire \bit_sel[22] ;
 wire \bit_sel[23] ;
 wire \bit_sel[24] ;
 wire \bit_sel[25] ;
 wire \bit_sel[26] ;
 wire \bit_sel[27] ;
 wire \bit_sel[28] ;
 wire \bit_sel[29] ;
 wire \bit_sel[2] ;
 wire \bit_sel[30] ;
 wire \bit_sel[31] ;
 wire \bit_sel[32] ;
 wire \bit_sel[33] ;
 wire \bit_sel[34] ;
 wire \bit_sel[35] ;
 wire \bit_sel[36] ;
 wire \bit_sel[37] ;
 wire \bit_sel[38] ;
 wire \bit_sel[39] ;
 wire \bit_sel[3] ;
 wire \bit_sel[40] ;
 wire \bit_sel[41] ;
 wire \bit_sel[42] ;
 wire \bit_sel[43] ;
 wire \bit_sel[44] ;
 wire \bit_sel[45] ;
 wire \bit_sel[46] ;
 wire \bit_sel[47] ;
 wire \bit_sel[48] ;
 wire \bit_sel[49] ;
 wire \bit_sel[4] ;
 wire \bit_sel[50] ;
 wire \bit_sel[51] ;
 wire \bit_sel[52] ;
 wire \bit_sel[53] ;
 wire \bit_sel[54] ;
 wire \bit_sel[55] ;
 wire \bit_sel[56] ;
 wire \bit_sel[57] ;
 wire \bit_sel[58] ;
 wire \bit_sel[59] ;
 wire \bit_sel[5] ;
 wire \bit_sel[60] ;
 wire \bit_sel[61] ;
 wire \bit_sel[62] ;
 wire \bit_sel[63] ;
 wire \bit_sel[6] ;
 wire \bit_sel[7] ;
 wire \bit_sel[8] ;
 wire \bit_sel[9] ;
 wire \bit_sel_reg[0] ;
 wire \bit_sel_reg[10] ;
 wire \bit_sel_reg[11] ;
 wire \bit_sel_reg[12] ;
 wire \bit_sel_reg[13] ;
 wire \bit_sel_reg[14] ;
 wire \bit_sel_reg[15] ;
 wire \bit_sel_reg[16] ;
 wire \bit_sel_reg[17] ;
 wire \bit_sel_reg[18] ;
 wire \bit_sel_reg[19] ;
 wire \bit_sel_reg[1] ;
 wire \bit_sel_reg[20] ;
 wire \bit_sel_reg[21] ;
 wire \bit_sel_reg[22] ;
 wire \bit_sel_reg[23] ;
 wire \bit_sel_reg[24] ;
 wire \bit_sel_reg[25] ;
 wire \bit_sel_reg[26] ;
 wire \bit_sel_reg[27] ;
 wire \bit_sel_reg[28] ;
 wire \bit_sel_reg[29] ;
 wire \bit_sel_reg[2] ;
 wire \bit_sel_reg[30] ;
 wire \bit_sel_reg[31] ;
 wire \bit_sel_reg[32] ;
 wire \bit_sel_reg[33] ;
 wire \bit_sel_reg[34] ;
 wire \bit_sel_reg[35] ;
 wire \bit_sel_reg[36] ;
 wire \bit_sel_reg[37] ;
 wire \bit_sel_reg[38] ;
 wire \bit_sel_reg[39] ;
 wire \bit_sel_reg[3] ;
 wire \bit_sel_reg[40] ;
 wire \bit_sel_reg[41] ;
 wire \bit_sel_reg[42] ;
 wire \bit_sel_reg[43] ;
 wire \bit_sel_reg[44] ;
 wire \bit_sel_reg[45] ;
 wire \bit_sel_reg[46] ;
 wire \bit_sel_reg[47] ;
 wire \bit_sel_reg[48] ;
 wire \bit_sel_reg[49] ;
 wire \bit_sel_reg[4] ;
 wire \bit_sel_reg[50] ;
 wire \bit_sel_reg[51] ;
 wire \bit_sel_reg[52] ;
 wire \bit_sel_reg[53] ;
 wire \bit_sel_reg[54] ;
 wire \bit_sel_reg[55] ;
 wire \bit_sel_reg[56] ;
 wire \bit_sel_reg[57] ;
 wire \bit_sel_reg[58] ;
 wire \bit_sel_reg[59] ;
 wire \bit_sel_reg[5] ;
 wire \bit_sel_reg[60] ;
 wire \bit_sel_reg[61] ;
 wire \bit_sel_reg[62] ;
 wire \bit_sel_reg[63] ;
 wire \bit_sel_reg[6] ;
 wire \bit_sel_reg[7] ;
 wire \bit_sel_reg[8] ;
 wire \bit_sel_reg[9] ;
 wire \col_prog_n[0] ;
 wire \col_prog_n[100] ;
 wire \col_prog_n[101] ;
 wire \col_prog_n[102] ;
 wire \col_prog_n[103] ;
 wire \col_prog_n[104] ;
 wire \col_prog_n[105] ;
 wire \col_prog_n[106] ;
 wire \col_prog_n[107] ;
 wire \col_prog_n[108] ;
 wire \col_prog_n[109] ;
 wire \col_prog_n[10] ;
 wire \col_prog_n[110] ;
 wire \col_prog_n[111] ;
 wire \col_prog_n[112] ;
 wire \col_prog_n[113] ;
 wire \col_prog_n[114] ;
 wire \col_prog_n[115] ;
 wire \col_prog_n[116] ;
 wire \col_prog_n[117] ;
 wire \col_prog_n[118] ;
 wire \col_prog_n[119] ;
 wire \col_prog_n[11] ;
 wire \col_prog_n[120] ;
 wire \col_prog_n[121] ;
 wire \col_prog_n[122] ;
 wire \col_prog_n[123] ;
 wire \col_prog_n[124] ;
 wire \col_prog_n[125] ;
 wire \col_prog_n[126] ;
 wire \col_prog_n[127] ;
 wire \col_prog_n[128] ;
 wire \col_prog_n[129] ;
 wire \col_prog_n[12] ;
 wire \col_prog_n[130] ;
 wire \col_prog_n[131] ;
 wire \col_prog_n[132] ;
 wire \col_prog_n[133] ;
 wire \col_prog_n[134] ;
 wire \col_prog_n[135] ;
 wire \col_prog_n[136] ;
 wire \col_prog_n[137] ;
 wire \col_prog_n[138] ;
 wire \col_prog_n[139] ;
 wire \col_prog_n[13] ;
 wire \col_prog_n[140] ;
 wire \col_prog_n[141] ;
 wire \col_prog_n[142] ;
 wire \col_prog_n[143] ;
 wire \col_prog_n[144] ;
 wire \col_prog_n[145] ;
 wire \col_prog_n[146] ;
 wire \col_prog_n[147] ;
 wire \col_prog_n[148] ;
 wire \col_prog_n[149] ;
 wire \col_prog_n[14] ;
 wire \col_prog_n[150] ;
 wire \col_prog_n[151] ;
 wire \col_prog_n[152] ;
 wire \col_prog_n[153] ;
 wire \col_prog_n[154] ;
 wire \col_prog_n[155] ;
 wire \col_prog_n[156] ;
 wire \col_prog_n[157] ;
 wire \col_prog_n[158] ;
 wire \col_prog_n[159] ;
 wire \col_prog_n[15] ;
 wire \col_prog_n[160] ;
 wire \col_prog_n[161] ;
 wire \col_prog_n[162] ;
 wire \col_prog_n[163] ;
 wire \col_prog_n[164] ;
 wire \col_prog_n[165] ;
 wire \col_prog_n[166] ;
 wire \col_prog_n[167] ;
 wire \col_prog_n[168] ;
 wire \col_prog_n[169] ;
 wire \col_prog_n[16] ;
 wire \col_prog_n[170] ;
 wire \col_prog_n[171] ;
 wire \col_prog_n[172] ;
 wire \col_prog_n[173] ;
 wire \col_prog_n[174] ;
 wire \col_prog_n[175] ;
 wire \col_prog_n[176] ;
 wire \col_prog_n[177] ;
 wire \col_prog_n[178] ;
 wire \col_prog_n[179] ;
 wire \col_prog_n[17] ;
 wire \col_prog_n[180] ;
 wire \col_prog_n[181] ;
 wire \col_prog_n[182] ;
 wire \col_prog_n[183] ;
 wire \col_prog_n[184] ;
 wire \col_prog_n[185] ;
 wire \col_prog_n[186] ;
 wire \col_prog_n[187] ;
 wire \col_prog_n[188] ;
 wire \col_prog_n[189] ;
 wire \col_prog_n[18] ;
 wire \col_prog_n[190] ;
 wire \col_prog_n[191] ;
 wire \col_prog_n[192] ;
 wire \col_prog_n[193] ;
 wire \col_prog_n[194] ;
 wire \col_prog_n[195] ;
 wire \col_prog_n[196] ;
 wire \col_prog_n[197] ;
 wire \col_prog_n[198] ;
 wire \col_prog_n[199] ;
 wire \col_prog_n[19] ;
 wire \col_prog_n[1] ;
 wire \col_prog_n[200] ;
 wire \col_prog_n[201] ;
 wire \col_prog_n[202] ;
 wire \col_prog_n[203] ;
 wire \col_prog_n[204] ;
 wire \col_prog_n[205] ;
 wire \col_prog_n[206] ;
 wire \col_prog_n[207] ;
 wire \col_prog_n[208] ;
 wire \col_prog_n[209] ;
 wire \col_prog_n[20] ;
 wire \col_prog_n[210] ;
 wire \col_prog_n[211] ;
 wire \col_prog_n[212] ;
 wire \col_prog_n[213] ;
 wire \col_prog_n[214] ;
 wire \col_prog_n[215] ;
 wire \col_prog_n[216] ;
 wire \col_prog_n[217] ;
 wire \col_prog_n[218] ;
 wire \col_prog_n[219] ;
 wire \col_prog_n[21] ;
 wire \col_prog_n[220] ;
 wire \col_prog_n[221] ;
 wire \col_prog_n[222] ;
 wire \col_prog_n[223] ;
 wire \col_prog_n[224] ;
 wire \col_prog_n[225] ;
 wire \col_prog_n[226] ;
 wire \col_prog_n[227] ;
 wire \col_prog_n[228] ;
 wire \col_prog_n[229] ;
 wire \col_prog_n[22] ;
 wire \col_prog_n[230] ;
 wire \col_prog_n[231] ;
 wire \col_prog_n[232] ;
 wire \col_prog_n[233] ;
 wire \col_prog_n[234] ;
 wire \col_prog_n[235] ;
 wire \col_prog_n[236] ;
 wire \col_prog_n[237] ;
 wire \col_prog_n[238] ;
 wire \col_prog_n[239] ;
 wire \col_prog_n[23] ;
 wire \col_prog_n[240] ;
 wire \col_prog_n[241] ;
 wire \col_prog_n[242] ;
 wire \col_prog_n[243] ;
 wire \col_prog_n[244] ;
 wire \col_prog_n[245] ;
 wire \col_prog_n[246] ;
 wire \col_prog_n[247] ;
 wire \col_prog_n[248] ;
 wire \col_prog_n[249] ;
 wire \col_prog_n[24] ;
 wire \col_prog_n[250] ;
 wire \col_prog_n[251] ;
 wire \col_prog_n[252] ;
 wire \col_prog_n[253] ;
 wire \col_prog_n[254] ;
 wire \col_prog_n[255] ;
 wire \col_prog_n[256] ;
 wire \col_prog_n[257] ;
 wire \col_prog_n[258] ;
 wire \col_prog_n[259] ;
 wire \col_prog_n[25] ;
 wire \col_prog_n[260] ;
 wire \col_prog_n[261] ;
 wire \col_prog_n[262] ;
 wire \col_prog_n[263] ;
 wire \col_prog_n[264] ;
 wire \col_prog_n[265] ;
 wire \col_prog_n[266] ;
 wire \col_prog_n[267] ;
 wire \col_prog_n[268] ;
 wire \col_prog_n[269] ;
 wire \col_prog_n[26] ;
 wire \col_prog_n[270] ;
 wire \col_prog_n[271] ;
 wire \col_prog_n[272] ;
 wire \col_prog_n[273] ;
 wire \col_prog_n[274] ;
 wire \col_prog_n[275] ;
 wire \col_prog_n[276] ;
 wire \col_prog_n[277] ;
 wire \col_prog_n[278] ;
 wire \col_prog_n[279] ;
 wire \col_prog_n[27] ;
 wire \col_prog_n[280] ;
 wire \col_prog_n[281] ;
 wire \col_prog_n[282] ;
 wire \col_prog_n[283] ;
 wire \col_prog_n[284] ;
 wire \col_prog_n[285] ;
 wire \col_prog_n[286] ;
 wire \col_prog_n[287] ;
 wire \col_prog_n[288] ;
 wire \col_prog_n[289] ;
 wire \col_prog_n[28] ;
 wire \col_prog_n[290] ;
 wire \col_prog_n[291] ;
 wire \col_prog_n[292] ;
 wire \col_prog_n[293] ;
 wire \col_prog_n[294] ;
 wire \col_prog_n[295] ;
 wire \col_prog_n[296] ;
 wire \col_prog_n[297] ;
 wire \col_prog_n[298] ;
 wire \col_prog_n[299] ;
 wire \col_prog_n[29] ;
 wire \col_prog_n[2] ;
 wire \col_prog_n[300] ;
 wire \col_prog_n[301] ;
 wire \col_prog_n[302] ;
 wire \col_prog_n[303] ;
 wire \col_prog_n[304] ;
 wire \col_prog_n[305] ;
 wire \col_prog_n[306] ;
 wire \col_prog_n[307] ;
 wire \col_prog_n[308] ;
 wire \col_prog_n[309] ;
 wire \col_prog_n[30] ;
 wire \col_prog_n[310] ;
 wire \col_prog_n[311] ;
 wire \col_prog_n[312] ;
 wire \col_prog_n[313] ;
 wire \col_prog_n[314] ;
 wire \col_prog_n[315] ;
 wire \col_prog_n[316] ;
 wire \col_prog_n[317] ;
 wire \col_prog_n[318] ;
 wire \col_prog_n[319] ;
 wire \col_prog_n[31] ;
 wire \col_prog_n[320] ;
 wire \col_prog_n[321] ;
 wire \col_prog_n[322] ;
 wire \col_prog_n[323] ;
 wire \col_prog_n[324] ;
 wire \col_prog_n[325] ;
 wire \col_prog_n[326] ;
 wire \col_prog_n[327] ;
 wire \col_prog_n[328] ;
 wire \col_prog_n[329] ;
 wire \col_prog_n[32] ;
 wire \col_prog_n[330] ;
 wire \col_prog_n[331] ;
 wire \col_prog_n[332] ;
 wire \col_prog_n[333] ;
 wire \col_prog_n[334] ;
 wire \col_prog_n[335] ;
 wire \col_prog_n[336] ;
 wire \col_prog_n[337] ;
 wire \col_prog_n[338] ;
 wire \col_prog_n[339] ;
 wire \col_prog_n[33] ;
 wire \col_prog_n[340] ;
 wire \col_prog_n[341] ;
 wire \col_prog_n[342] ;
 wire \col_prog_n[343] ;
 wire \col_prog_n[344] ;
 wire \col_prog_n[345] ;
 wire \col_prog_n[346] ;
 wire \col_prog_n[347] ;
 wire \col_prog_n[348] ;
 wire \col_prog_n[349] ;
 wire \col_prog_n[34] ;
 wire \col_prog_n[350] ;
 wire \col_prog_n[351] ;
 wire \col_prog_n[352] ;
 wire \col_prog_n[353] ;
 wire \col_prog_n[354] ;
 wire \col_prog_n[355] ;
 wire \col_prog_n[356] ;
 wire \col_prog_n[357] ;
 wire \col_prog_n[358] ;
 wire \col_prog_n[359] ;
 wire \col_prog_n[35] ;
 wire \col_prog_n[360] ;
 wire \col_prog_n[361] ;
 wire \col_prog_n[362] ;
 wire \col_prog_n[363] ;
 wire \col_prog_n[364] ;
 wire \col_prog_n[365] ;
 wire \col_prog_n[366] ;
 wire \col_prog_n[367] ;
 wire \col_prog_n[368] ;
 wire \col_prog_n[369] ;
 wire \col_prog_n[36] ;
 wire \col_prog_n[370] ;
 wire \col_prog_n[371] ;
 wire \col_prog_n[372] ;
 wire \col_prog_n[373] ;
 wire \col_prog_n[374] ;
 wire \col_prog_n[375] ;
 wire \col_prog_n[376] ;
 wire \col_prog_n[377] ;
 wire \col_prog_n[378] ;
 wire \col_prog_n[379] ;
 wire \col_prog_n[37] ;
 wire \col_prog_n[380] ;
 wire \col_prog_n[381] ;
 wire \col_prog_n[382] ;
 wire \col_prog_n[383] ;
 wire \col_prog_n[384] ;
 wire \col_prog_n[385] ;
 wire \col_prog_n[386] ;
 wire \col_prog_n[387] ;
 wire \col_prog_n[388] ;
 wire \col_prog_n[389] ;
 wire \col_prog_n[38] ;
 wire \col_prog_n[390] ;
 wire \col_prog_n[391] ;
 wire \col_prog_n[392] ;
 wire \col_prog_n[393] ;
 wire \col_prog_n[394] ;
 wire \col_prog_n[395] ;
 wire \col_prog_n[396] ;
 wire \col_prog_n[397] ;
 wire \col_prog_n[398] ;
 wire \col_prog_n[399] ;
 wire \col_prog_n[39] ;
 wire \col_prog_n[3] ;
 wire \col_prog_n[400] ;
 wire \col_prog_n[401] ;
 wire \col_prog_n[402] ;
 wire \col_prog_n[403] ;
 wire \col_prog_n[404] ;
 wire \col_prog_n[405] ;
 wire \col_prog_n[406] ;
 wire \col_prog_n[407] ;
 wire \col_prog_n[408] ;
 wire \col_prog_n[409] ;
 wire \col_prog_n[40] ;
 wire \col_prog_n[410] ;
 wire \col_prog_n[411] ;
 wire \col_prog_n[412] ;
 wire \col_prog_n[413] ;
 wire \col_prog_n[414] ;
 wire \col_prog_n[415] ;
 wire \col_prog_n[416] ;
 wire \col_prog_n[417] ;
 wire \col_prog_n[418] ;
 wire \col_prog_n[419] ;
 wire \col_prog_n[41] ;
 wire \col_prog_n[420] ;
 wire \col_prog_n[421] ;
 wire \col_prog_n[422] ;
 wire \col_prog_n[423] ;
 wire \col_prog_n[424] ;
 wire \col_prog_n[425] ;
 wire \col_prog_n[426] ;
 wire \col_prog_n[427] ;
 wire \col_prog_n[428] ;
 wire \col_prog_n[429] ;
 wire \col_prog_n[42] ;
 wire \col_prog_n[430] ;
 wire \col_prog_n[431] ;
 wire \col_prog_n[432] ;
 wire \col_prog_n[433] ;
 wire \col_prog_n[434] ;
 wire \col_prog_n[435] ;
 wire \col_prog_n[436] ;
 wire \col_prog_n[437] ;
 wire \col_prog_n[438] ;
 wire \col_prog_n[439] ;
 wire \col_prog_n[43] ;
 wire \col_prog_n[440] ;
 wire \col_prog_n[441] ;
 wire \col_prog_n[442] ;
 wire \col_prog_n[443] ;
 wire \col_prog_n[444] ;
 wire \col_prog_n[445] ;
 wire \col_prog_n[446] ;
 wire \col_prog_n[447] ;
 wire \col_prog_n[448] ;
 wire \col_prog_n[449] ;
 wire \col_prog_n[44] ;
 wire \col_prog_n[450] ;
 wire \col_prog_n[451] ;
 wire \col_prog_n[452] ;
 wire \col_prog_n[453] ;
 wire \col_prog_n[454] ;
 wire \col_prog_n[455] ;
 wire \col_prog_n[456] ;
 wire \col_prog_n[457] ;
 wire \col_prog_n[458] ;
 wire \col_prog_n[459] ;
 wire \col_prog_n[45] ;
 wire \col_prog_n[460] ;
 wire \col_prog_n[461] ;
 wire \col_prog_n[462] ;
 wire \col_prog_n[463] ;
 wire \col_prog_n[464] ;
 wire \col_prog_n[465] ;
 wire \col_prog_n[466] ;
 wire \col_prog_n[467] ;
 wire \col_prog_n[468] ;
 wire \col_prog_n[469] ;
 wire \col_prog_n[46] ;
 wire \col_prog_n[470] ;
 wire \col_prog_n[471] ;
 wire \col_prog_n[472] ;
 wire \col_prog_n[473] ;
 wire \col_prog_n[474] ;
 wire \col_prog_n[475] ;
 wire \col_prog_n[476] ;
 wire \col_prog_n[477] ;
 wire \col_prog_n[478] ;
 wire \col_prog_n[479] ;
 wire \col_prog_n[47] ;
 wire \col_prog_n[480] ;
 wire \col_prog_n[481] ;
 wire \col_prog_n[482] ;
 wire \col_prog_n[483] ;
 wire \col_prog_n[484] ;
 wire \col_prog_n[485] ;
 wire \col_prog_n[486] ;
 wire \col_prog_n[487] ;
 wire \col_prog_n[488] ;
 wire \col_prog_n[489] ;
 wire \col_prog_n[48] ;
 wire \col_prog_n[490] ;
 wire \col_prog_n[491] ;
 wire \col_prog_n[492] ;
 wire \col_prog_n[493] ;
 wire \col_prog_n[494] ;
 wire \col_prog_n[495] ;
 wire \col_prog_n[496] ;
 wire \col_prog_n[497] ;
 wire \col_prog_n[498] ;
 wire \col_prog_n[499] ;
 wire \col_prog_n[49] ;
 wire \col_prog_n[4] ;
 wire \col_prog_n[500] ;
 wire \col_prog_n[501] ;
 wire \col_prog_n[502] ;
 wire \col_prog_n[503] ;
 wire \col_prog_n[504] ;
 wire \col_prog_n[505] ;
 wire \col_prog_n[506] ;
 wire \col_prog_n[507] ;
 wire \col_prog_n[508] ;
 wire \col_prog_n[509] ;
 wire \col_prog_n[50] ;
 wire \col_prog_n[510] ;
 wire \col_prog_n[511] ;
 wire \col_prog_n[51] ;
 wire \col_prog_n[52] ;
 wire \col_prog_n[53] ;
 wire \col_prog_n[54] ;
 wire \col_prog_n[55] ;
 wire \col_prog_n[56] ;
 wire \col_prog_n[57] ;
 wire \col_prog_n[58] ;
 wire \col_prog_n[59] ;
 wire \col_prog_n[5] ;
 wire \col_prog_n[60] ;
 wire \col_prog_n[61] ;
 wire \col_prog_n[62] ;
 wire \col_prog_n[63] ;
 wire \col_prog_n[64] ;
 wire \col_prog_n[65] ;
 wire \col_prog_n[66] ;
 wire \col_prog_n[67] ;
 wire \col_prog_n[68] ;
 wire \col_prog_n[69] ;
 wire \col_prog_n[6] ;
 wire \col_prog_n[70] ;
 wire \col_prog_n[71] ;
 wire \col_prog_n[72] ;
 wire \col_prog_n[73] ;
 wire \col_prog_n[74] ;
 wire \col_prog_n[75] ;
 wire \col_prog_n[76] ;
 wire \col_prog_n[77] ;
 wire \col_prog_n[78] ;
 wire \col_prog_n[79] ;
 wire \col_prog_n[7] ;
 wire \col_prog_n[80] ;
 wire \col_prog_n[81] ;
 wire \col_prog_n[82] ;
 wire \col_prog_n[83] ;
 wire \col_prog_n[84] ;
 wire \col_prog_n[85] ;
 wire \col_prog_n[86] ;
 wire \col_prog_n[87] ;
 wire \col_prog_n[88] ;
 wire \col_prog_n[89] ;
 wire \col_prog_n[8] ;
 wire \col_prog_n[90] ;
 wire \col_prog_n[91] ;
 wire \col_prog_n[92] ;
 wire \col_prog_n[93] ;
 wire \col_prog_n[94] ;
 wire \col_prog_n[95] ;
 wire \col_prog_n[96] ;
 wire \col_prog_n[97] ;
 wire \col_prog_n[98] ;
 wire \col_prog_n[99] ;
 wire \col_prog_n[9] ;
 wire \col_prog_n_reg[0] ;
 wire \col_prog_n_reg[100] ;
 wire \col_prog_n_reg[101] ;
 wire \col_prog_n_reg[102] ;
 wire \col_prog_n_reg[103] ;
 wire \col_prog_n_reg[104] ;
 wire \col_prog_n_reg[105] ;
 wire \col_prog_n_reg[106] ;
 wire \col_prog_n_reg[107] ;
 wire \col_prog_n_reg[108] ;
 wire \col_prog_n_reg[109] ;
 wire \col_prog_n_reg[10] ;
 wire \col_prog_n_reg[110] ;
 wire \col_prog_n_reg[111] ;
 wire \col_prog_n_reg[112] ;
 wire \col_prog_n_reg[113] ;
 wire \col_prog_n_reg[114] ;
 wire \col_prog_n_reg[115] ;
 wire \col_prog_n_reg[116] ;
 wire \col_prog_n_reg[117] ;
 wire \col_prog_n_reg[118] ;
 wire \col_prog_n_reg[119] ;
 wire \col_prog_n_reg[11] ;
 wire \col_prog_n_reg[120] ;
 wire \col_prog_n_reg[121] ;
 wire \col_prog_n_reg[122] ;
 wire \col_prog_n_reg[123] ;
 wire \col_prog_n_reg[124] ;
 wire \col_prog_n_reg[125] ;
 wire \col_prog_n_reg[126] ;
 wire \col_prog_n_reg[127] ;
 wire \col_prog_n_reg[128] ;
 wire \col_prog_n_reg[129] ;
 wire \col_prog_n_reg[12] ;
 wire \col_prog_n_reg[130] ;
 wire \col_prog_n_reg[131] ;
 wire \col_prog_n_reg[132] ;
 wire \col_prog_n_reg[133] ;
 wire \col_prog_n_reg[134] ;
 wire \col_prog_n_reg[135] ;
 wire \col_prog_n_reg[136] ;
 wire \col_prog_n_reg[137] ;
 wire \col_prog_n_reg[138] ;
 wire \col_prog_n_reg[139] ;
 wire \col_prog_n_reg[13] ;
 wire \col_prog_n_reg[140] ;
 wire \col_prog_n_reg[141] ;
 wire \col_prog_n_reg[142] ;
 wire \col_prog_n_reg[143] ;
 wire \col_prog_n_reg[144] ;
 wire \col_prog_n_reg[145] ;
 wire \col_prog_n_reg[146] ;
 wire \col_prog_n_reg[147] ;
 wire \col_prog_n_reg[148] ;
 wire \col_prog_n_reg[149] ;
 wire \col_prog_n_reg[14] ;
 wire \col_prog_n_reg[150] ;
 wire \col_prog_n_reg[151] ;
 wire \col_prog_n_reg[152] ;
 wire \col_prog_n_reg[153] ;
 wire \col_prog_n_reg[154] ;
 wire \col_prog_n_reg[155] ;
 wire \col_prog_n_reg[156] ;
 wire \col_prog_n_reg[157] ;
 wire \col_prog_n_reg[158] ;
 wire \col_prog_n_reg[159] ;
 wire \col_prog_n_reg[15] ;
 wire \col_prog_n_reg[160] ;
 wire \col_prog_n_reg[161] ;
 wire \col_prog_n_reg[162] ;
 wire \col_prog_n_reg[163] ;
 wire \col_prog_n_reg[164] ;
 wire \col_prog_n_reg[165] ;
 wire \col_prog_n_reg[166] ;
 wire \col_prog_n_reg[167] ;
 wire \col_prog_n_reg[168] ;
 wire \col_prog_n_reg[169] ;
 wire \col_prog_n_reg[16] ;
 wire \col_prog_n_reg[170] ;
 wire \col_prog_n_reg[171] ;
 wire \col_prog_n_reg[172] ;
 wire \col_prog_n_reg[173] ;
 wire \col_prog_n_reg[174] ;
 wire \col_prog_n_reg[175] ;
 wire \col_prog_n_reg[176] ;
 wire \col_prog_n_reg[177] ;
 wire \col_prog_n_reg[178] ;
 wire \col_prog_n_reg[179] ;
 wire \col_prog_n_reg[17] ;
 wire \col_prog_n_reg[180] ;
 wire \col_prog_n_reg[181] ;
 wire \col_prog_n_reg[182] ;
 wire \col_prog_n_reg[183] ;
 wire \col_prog_n_reg[184] ;
 wire \col_prog_n_reg[185] ;
 wire \col_prog_n_reg[186] ;
 wire \col_prog_n_reg[187] ;
 wire \col_prog_n_reg[188] ;
 wire \col_prog_n_reg[189] ;
 wire \col_prog_n_reg[18] ;
 wire \col_prog_n_reg[190] ;
 wire \col_prog_n_reg[191] ;
 wire \col_prog_n_reg[192] ;
 wire \col_prog_n_reg[193] ;
 wire \col_prog_n_reg[194] ;
 wire \col_prog_n_reg[195] ;
 wire \col_prog_n_reg[196] ;
 wire \col_prog_n_reg[197] ;
 wire \col_prog_n_reg[198] ;
 wire \col_prog_n_reg[199] ;
 wire \col_prog_n_reg[19] ;
 wire \col_prog_n_reg[1] ;
 wire \col_prog_n_reg[200] ;
 wire \col_prog_n_reg[201] ;
 wire \col_prog_n_reg[202] ;
 wire \col_prog_n_reg[203] ;
 wire \col_prog_n_reg[204] ;
 wire \col_prog_n_reg[205] ;
 wire \col_prog_n_reg[206] ;
 wire \col_prog_n_reg[207] ;
 wire \col_prog_n_reg[208] ;
 wire \col_prog_n_reg[209] ;
 wire \col_prog_n_reg[20] ;
 wire \col_prog_n_reg[210] ;
 wire \col_prog_n_reg[211] ;
 wire \col_prog_n_reg[212] ;
 wire \col_prog_n_reg[213] ;
 wire \col_prog_n_reg[214] ;
 wire \col_prog_n_reg[215] ;
 wire \col_prog_n_reg[216] ;
 wire \col_prog_n_reg[217] ;
 wire \col_prog_n_reg[218] ;
 wire \col_prog_n_reg[219] ;
 wire \col_prog_n_reg[21] ;
 wire \col_prog_n_reg[220] ;
 wire \col_prog_n_reg[221] ;
 wire \col_prog_n_reg[222] ;
 wire \col_prog_n_reg[223] ;
 wire \col_prog_n_reg[224] ;
 wire \col_prog_n_reg[225] ;
 wire \col_prog_n_reg[226] ;
 wire \col_prog_n_reg[227] ;
 wire \col_prog_n_reg[228] ;
 wire \col_prog_n_reg[229] ;
 wire \col_prog_n_reg[22] ;
 wire \col_prog_n_reg[230] ;
 wire \col_prog_n_reg[231] ;
 wire \col_prog_n_reg[232] ;
 wire \col_prog_n_reg[233] ;
 wire \col_prog_n_reg[234] ;
 wire \col_prog_n_reg[235] ;
 wire \col_prog_n_reg[236] ;
 wire \col_prog_n_reg[237] ;
 wire \col_prog_n_reg[238] ;
 wire \col_prog_n_reg[239] ;
 wire \col_prog_n_reg[23] ;
 wire \col_prog_n_reg[240] ;
 wire \col_prog_n_reg[241] ;
 wire \col_prog_n_reg[242] ;
 wire \col_prog_n_reg[243] ;
 wire \col_prog_n_reg[244] ;
 wire \col_prog_n_reg[245] ;
 wire \col_prog_n_reg[246] ;
 wire \col_prog_n_reg[247] ;
 wire \col_prog_n_reg[248] ;
 wire \col_prog_n_reg[249] ;
 wire \col_prog_n_reg[24] ;
 wire \col_prog_n_reg[250] ;
 wire \col_prog_n_reg[251] ;
 wire \col_prog_n_reg[252] ;
 wire \col_prog_n_reg[253] ;
 wire \col_prog_n_reg[254] ;
 wire \col_prog_n_reg[255] ;
 wire \col_prog_n_reg[256] ;
 wire \col_prog_n_reg[257] ;
 wire \col_prog_n_reg[258] ;
 wire \col_prog_n_reg[259] ;
 wire \col_prog_n_reg[25] ;
 wire \col_prog_n_reg[260] ;
 wire \col_prog_n_reg[261] ;
 wire \col_prog_n_reg[262] ;
 wire \col_prog_n_reg[263] ;
 wire \col_prog_n_reg[264] ;
 wire \col_prog_n_reg[265] ;
 wire \col_prog_n_reg[266] ;
 wire \col_prog_n_reg[267] ;
 wire \col_prog_n_reg[268] ;
 wire \col_prog_n_reg[269] ;
 wire \col_prog_n_reg[26] ;
 wire \col_prog_n_reg[270] ;
 wire \col_prog_n_reg[271] ;
 wire \col_prog_n_reg[272] ;
 wire \col_prog_n_reg[273] ;
 wire \col_prog_n_reg[274] ;
 wire \col_prog_n_reg[275] ;
 wire \col_prog_n_reg[276] ;
 wire \col_prog_n_reg[277] ;
 wire \col_prog_n_reg[278] ;
 wire \col_prog_n_reg[279] ;
 wire \col_prog_n_reg[27] ;
 wire \col_prog_n_reg[280] ;
 wire \col_prog_n_reg[281] ;
 wire \col_prog_n_reg[282] ;
 wire \col_prog_n_reg[283] ;
 wire \col_prog_n_reg[284] ;
 wire \col_prog_n_reg[285] ;
 wire \col_prog_n_reg[286] ;
 wire \col_prog_n_reg[287] ;
 wire \col_prog_n_reg[288] ;
 wire \col_prog_n_reg[289] ;
 wire \col_prog_n_reg[28] ;
 wire \col_prog_n_reg[290] ;
 wire \col_prog_n_reg[291] ;
 wire \col_prog_n_reg[292] ;
 wire \col_prog_n_reg[293] ;
 wire \col_prog_n_reg[294] ;
 wire \col_prog_n_reg[295] ;
 wire \col_prog_n_reg[296] ;
 wire \col_prog_n_reg[297] ;
 wire \col_prog_n_reg[298] ;
 wire \col_prog_n_reg[299] ;
 wire \col_prog_n_reg[29] ;
 wire \col_prog_n_reg[2] ;
 wire \col_prog_n_reg[300] ;
 wire \col_prog_n_reg[301] ;
 wire \col_prog_n_reg[302] ;
 wire \col_prog_n_reg[303] ;
 wire \col_prog_n_reg[304] ;
 wire \col_prog_n_reg[305] ;
 wire \col_prog_n_reg[306] ;
 wire \col_prog_n_reg[307] ;
 wire \col_prog_n_reg[308] ;
 wire \col_prog_n_reg[309] ;
 wire \col_prog_n_reg[30] ;
 wire \col_prog_n_reg[310] ;
 wire \col_prog_n_reg[311] ;
 wire \col_prog_n_reg[312] ;
 wire \col_prog_n_reg[313] ;
 wire \col_prog_n_reg[314] ;
 wire \col_prog_n_reg[315] ;
 wire \col_prog_n_reg[316] ;
 wire \col_prog_n_reg[317] ;
 wire \col_prog_n_reg[318] ;
 wire \col_prog_n_reg[319] ;
 wire \col_prog_n_reg[31] ;
 wire \col_prog_n_reg[320] ;
 wire \col_prog_n_reg[321] ;
 wire \col_prog_n_reg[322] ;
 wire \col_prog_n_reg[323] ;
 wire \col_prog_n_reg[324] ;
 wire \col_prog_n_reg[325] ;
 wire \col_prog_n_reg[326] ;
 wire \col_prog_n_reg[327] ;
 wire \col_prog_n_reg[328] ;
 wire \col_prog_n_reg[329] ;
 wire \col_prog_n_reg[32] ;
 wire \col_prog_n_reg[330] ;
 wire \col_prog_n_reg[331] ;
 wire \col_prog_n_reg[332] ;
 wire \col_prog_n_reg[333] ;
 wire \col_prog_n_reg[334] ;
 wire \col_prog_n_reg[335] ;
 wire \col_prog_n_reg[336] ;
 wire \col_prog_n_reg[337] ;
 wire \col_prog_n_reg[338] ;
 wire \col_prog_n_reg[339] ;
 wire \col_prog_n_reg[33] ;
 wire \col_prog_n_reg[340] ;
 wire \col_prog_n_reg[341] ;
 wire \col_prog_n_reg[342] ;
 wire \col_prog_n_reg[343] ;
 wire \col_prog_n_reg[344] ;
 wire \col_prog_n_reg[345] ;
 wire \col_prog_n_reg[346] ;
 wire \col_prog_n_reg[347] ;
 wire \col_prog_n_reg[348] ;
 wire \col_prog_n_reg[349] ;
 wire \col_prog_n_reg[34] ;
 wire \col_prog_n_reg[350] ;
 wire \col_prog_n_reg[351] ;
 wire \col_prog_n_reg[352] ;
 wire \col_prog_n_reg[353] ;
 wire \col_prog_n_reg[354] ;
 wire \col_prog_n_reg[355] ;
 wire \col_prog_n_reg[356] ;
 wire \col_prog_n_reg[357] ;
 wire \col_prog_n_reg[358] ;
 wire \col_prog_n_reg[359] ;
 wire \col_prog_n_reg[35] ;
 wire \col_prog_n_reg[360] ;
 wire \col_prog_n_reg[361] ;
 wire \col_prog_n_reg[362] ;
 wire \col_prog_n_reg[363] ;
 wire \col_prog_n_reg[364] ;
 wire \col_prog_n_reg[365] ;
 wire \col_prog_n_reg[366] ;
 wire \col_prog_n_reg[367] ;
 wire \col_prog_n_reg[368] ;
 wire \col_prog_n_reg[369] ;
 wire \col_prog_n_reg[36] ;
 wire \col_prog_n_reg[370] ;
 wire \col_prog_n_reg[371] ;
 wire \col_prog_n_reg[372] ;
 wire \col_prog_n_reg[373] ;
 wire \col_prog_n_reg[374] ;
 wire \col_prog_n_reg[375] ;
 wire \col_prog_n_reg[376] ;
 wire \col_prog_n_reg[377] ;
 wire \col_prog_n_reg[378] ;
 wire \col_prog_n_reg[379] ;
 wire \col_prog_n_reg[37] ;
 wire \col_prog_n_reg[380] ;
 wire \col_prog_n_reg[381] ;
 wire \col_prog_n_reg[382] ;
 wire \col_prog_n_reg[383] ;
 wire \col_prog_n_reg[384] ;
 wire \col_prog_n_reg[385] ;
 wire \col_prog_n_reg[386] ;
 wire \col_prog_n_reg[387] ;
 wire \col_prog_n_reg[388] ;
 wire \col_prog_n_reg[389] ;
 wire \col_prog_n_reg[38] ;
 wire \col_prog_n_reg[390] ;
 wire \col_prog_n_reg[391] ;
 wire \col_prog_n_reg[392] ;
 wire \col_prog_n_reg[393] ;
 wire \col_prog_n_reg[394] ;
 wire \col_prog_n_reg[395] ;
 wire \col_prog_n_reg[396] ;
 wire \col_prog_n_reg[397] ;
 wire \col_prog_n_reg[398] ;
 wire \col_prog_n_reg[399] ;
 wire \col_prog_n_reg[39] ;
 wire \col_prog_n_reg[3] ;
 wire \col_prog_n_reg[400] ;
 wire \col_prog_n_reg[401] ;
 wire \col_prog_n_reg[402] ;
 wire \col_prog_n_reg[403] ;
 wire \col_prog_n_reg[404] ;
 wire \col_prog_n_reg[405] ;
 wire \col_prog_n_reg[406] ;
 wire \col_prog_n_reg[407] ;
 wire \col_prog_n_reg[408] ;
 wire \col_prog_n_reg[409] ;
 wire \col_prog_n_reg[40] ;
 wire \col_prog_n_reg[410] ;
 wire \col_prog_n_reg[411] ;
 wire \col_prog_n_reg[412] ;
 wire \col_prog_n_reg[413] ;
 wire \col_prog_n_reg[414] ;
 wire \col_prog_n_reg[415] ;
 wire \col_prog_n_reg[416] ;
 wire \col_prog_n_reg[417] ;
 wire \col_prog_n_reg[418] ;
 wire \col_prog_n_reg[419] ;
 wire \col_prog_n_reg[41] ;
 wire \col_prog_n_reg[420] ;
 wire \col_prog_n_reg[421] ;
 wire \col_prog_n_reg[422] ;
 wire \col_prog_n_reg[423] ;
 wire \col_prog_n_reg[424] ;
 wire \col_prog_n_reg[425] ;
 wire \col_prog_n_reg[426] ;
 wire \col_prog_n_reg[427] ;
 wire \col_prog_n_reg[428] ;
 wire \col_prog_n_reg[429] ;
 wire \col_prog_n_reg[42] ;
 wire \col_prog_n_reg[430] ;
 wire \col_prog_n_reg[431] ;
 wire \col_prog_n_reg[432] ;
 wire \col_prog_n_reg[433] ;
 wire \col_prog_n_reg[434] ;
 wire \col_prog_n_reg[435] ;
 wire \col_prog_n_reg[436] ;
 wire \col_prog_n_reg[437] ;
 wire \col_prog_n_reg[438] ;
 wire \col_prog_n_reg[439] ;
 wire \col_prog_n_reg[43] ;
 wire \col_prog_n_reg[440] ;
 wire \col_prog_n_reg[441] ;
 wire \col_prog_n_reg[442] ;
 wire \col_prog_n_reg[443] ;
 wire \col_prog_n_reg[444] ;
 wire \col_prog_n_reg[445] ;
 wire \col_prog_n_reg[446] ;
 wire \col_prog_n_reg[447] ;
 wire \col_prog_n_reg[448] ;
 wire \col_prog_n_reg[449] ;
 wire \col_prog_n_reg[44] ;
 wire \col_prog_n_reg[450] ;
 wire \col_prog_n_reg[451] ;
 wire \col_prog_n_reg[452] ;
 wire \col_prog_n_reg[453] ;
 wire \col_prog_n_reg[454] ;
 wire \col_prog_n_reg[455] ;
 wire \col_prog_n_reg[456] ;
 wire \col_prog_n_reg[457] ;
 wire \col_prog_n_reg[458] ;
 wire \col_prog_n_reg[459] ;
 wire \col_prog_n_reg[45] ;
 wire \col_prog_n_reg[460] ;
 wire \col_prog_n_reg[461] ;
 wire \col_prog_n_reg[462] ;
 wire \col_prog_n_reg[463] ;
 wire \col_prog_n_reg[464] ;
 wire \col_prog_n_reg[465] ;
 wire \col_prog_n_reg[466] ;
 wire \col_prog_n_reg[467] ;
 wire \col_prog_n_reg[468] ;
 wire \col_prog_n_reg[469] ;
 wire \col_prog_n_reg[46] ;
 wire \col_prog_n_reg[470] ;
 wire \col_prog_n_reg[471] ;
 wire \col_prog_n_reg[472] ;
 wire \col_prog_n_reg[473] ;
 wire \col_prog_n_reg[474] ;
 wire \col_prog_n_reg[475] ;
 wire \col_prog_n_reg[476] ;
 wire \col_prog_n_reg[477] ;
 wire \col_prog_n_reg[478] ;
 wire \col_prog_n_reg[479] ;
 wire \col_prog_n_reg[47] ;
 wire \col_prog_n_reg[480] ;
 wire \col_prog_n_reg[481] ;
 wire \col_prog_n_reg[482] ;
 wire \col_prog_n_reg[483] ;
 wire \col_prog_n_reg[484] ;
 wire \col_prog_n_reg[485] ;
 wire \col_prog_n_reg[486] ;
 wire \col_prog_n_reg[487] ;
 wire \col_prog_n_reg[488] ;
 wire \col_prog_n_reg[489] ;
 wire \col_prog_n_reg[48] ;
 wire \col_prog_n_reg[490] ;
 wire \col_prog_n_reg[491] ;
 wire \col_prog_n_reg[492] ;
 wire \col_prog_n_reg[493] ;
 wire \col_prog_n_reg[494] ;
 wire \col_prog_n_reg[495] ;
 wire \col_prog_n_reg[496] ;
 wire \col_prog_n_reg[497] ;
 wire \col_prog_n_reg[498] ;
 wire \col_prog_n_reg[499] ;
 wire \col_prog_n_reg[49] ;
 wire \col_prog_n_reg[4] ;
 wire \col_prog_n_reg[500] ;
 wire \col_prog_n_reg[501] ;
 wire \col_prog_n_reg[502] ;
 wire \col_prog_n_reg[503] ;
 wire \col_prog_n_reg[504] ;
 wire \col_prog_n_reg[505] ;
 wire \col_prog_n_reg[506] ;
 wire \col_prog_n_reg[507] ;
 wire \col_prog_n_reg[508] ;
 wire \col_prog_n_reg[509] ;
 wire \col_prog_n_reg[50] ;
 wire \col_prog_n_reg[510] ;
 wire \col_prog_n_reg[511] ;
 wire \col_prog_n_reg[51] ;
 wire \col_prog_n_reg[52] ;
 wire \col_prog_n_reg[53] ;
 wire \col_prog_n_reg[54] ;
 wire \col_prog_n_reg[55] ;
 wire \col_prog_n_reg[56] ;
 wire \col_prog_n_reg[57] ;
 wire \col_prog_n_reg[58] ;
 wire \col_prog_n_reg[59] ;
 wire \col_prog_n_reg[5] ;
 wire \col_prog_n_reg[60] ;
 wire \col_prog_n_reg[61] ;
 wire \col_prog_n_reg[62] ;
 wire \col_prog_n_reg[63] ;
 wire \col_prog_n_reg[64] ;
 wire \col_prog_n_reg[65] ;
 wire \col_prog_n_reg[66] ;
 wire \col_prog_n_reg[67] ;
 wire \col_prog_n_reg[68] ;
 wire \col_prog_n_reg[69] ;
 wire \col_prog_n_reg[6] ;
 wire \col_prog_n_reg[70] ;
 wire \col_prog_n_reg[71] ;
 wire \col_prog_n_reg[72] ;
 wire \col_prog_n_reg[73] ;
 wire \col_prog_n_reg[74] ;
 wire \col_prog_n_reg[75] ;
 wire \col_prog_n_reg[76] ;
 wire \col_prog_n_reg[77] ;
 wire \col_prog_n_reg[78] ;
 wire \col_prog_n_reg[79] ;
 wire \col_prog_n_reg[7] ;
 wire \col_prog_n_reg[80] ;
 wire \col_prog_n_reg[81] ;
 wire \col_prog_n_reg[82] ;
 wire \col_prog_n_reg[83] ;
 wire \col_prog_n_reg[84] ;
 wire \col_prog_n_reg[85] ;
 wire \col_prog_n_reg[86] ;
 wire \col_prog_n_reg[87] ;
 wire \col_prog_n_reg[88] ;
 wire \col_prog_n_reg[89] ;
 wire \col_prog_n_reg[8] ;
 wire \col_prog_n_reg[90] ;
 wire \col_prog_n_reg[91] ;
 wire \col_prog_n_reg[92] ;
 wire \col_prog_n_reg[93] ;
 wire \col_prog_n_reg[94] ;
 wire \col_prog_n_reg[95] ;
 wire \col_prog_n_reg[96] ;
 wire \col_prog_n_reg[97] ;
 wire \col_prog_n_reg[98] ;
 wire \col_prog_n_reg[99] ;
 wire \col_prog_n_reg[9] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \efuse_out[0] ;
 wire \efuse_out[100] ;
 wire \efuse_out[101] ;
 wire \efuse_out[102] ;
 wire \efuse_out[103] ;
 wire \efuse_out[104] ;
 wire \efuse_out[105] ;
 wire \efuse_out[106] ;
 wire \efuse_out[107] ;
 wire \efuse_out[108] ;
 wire \efuse_out[109] ;
 wire \efuse_out[10] ;
 wire \efuse_out[110] ;
 wire \efuse_out[111] ;
 wire \efuse_out[112] ;
 wire \efuse_out[113] ;
 wire \efuse_out[114] ;
 wire \efuse_out[115] ;
 wire \efuse_out[116] ;
 wire \efuse_out[117] ;
 wire \efuse_out[118] ;
 wire \efuse_out[119] ;
 wire \efuse_out[11] ;
 wire \efuse_out[120] ;
 wire \efuse_out[121] ;
 wire \efuse_out[122] ;
 wire \efuse_out[123] ;
 wire \efuse_out[124] ;
 wire \efuse_out[125] ;
 wire \efuse_out[126] ;
 wire \efuse_out[127] ;
 wire \efuse_out[128] ;
 wire \efuse_out[129] ;
 wire \efuse_out[12] ;
 wire \efuse_out[130] ;
 wire \efuse_out[131] ;
 wire \efuse_out[132] ;
 wire \efuse_out[133] ;
 wire \efuse_out[134] ;
 wire \efuse_out[135] ;
 wire \efuse_out[136] ;
 wire \efuse_out[137] ;
 wire \efuse_out[138] ;
 wire \efuse_out[139] ;
 wire \efuse_out[13] ;
 wire \efuse_out[140] ;
 wire \efuse_out[141] ;
 wire \efuse_out[142] ;
 wire \efuse_out[143] ;
 wire \efuse_out[144] ;
 wire \efuse_out[145] ;
 wire \efuse_out[146] ;
 wire \efuse_out[147] ;
 wire \efuse_out[148] ;
 wire \efuse_out[149] ;
 wire \efuse_out[14] ;
 wire \efuse_out[150] ;
 wire \efuse_out[151] ;
 wire \efuse_out[152] ;
 wire \efuse_out[153] ;
 wire \efuse_out[154] ;
 wire \efuse_out[155] ;
 wire \efuse_out[156] ;
 wire \efuse_out[157] ;
 wire \efuse_out[158] ;
 wire \efuse_out[159] ;
 wire \efuse_out[15] ;
 wire \efuse_out[160] ;
 wire \efuse_out[161] ;
 wire \efuse_out[162] ;
 wire \efuse_out[163] ;
 wire \efuse_out[164] ;
 wire \efuse_out[165] ;
 wire \efuse_out[166] ;
 wire \efuse_out[167] ;
 wire \efuse_out[168] ;
 wire \efuse_out[169] ;
 wire \efuse_out[16] ;
 wire \efuse_out[170] ;
 wire \efuse_out[171] ;
 wire \efuse_out[172] ;
 wire \efuse_out[173] ;
 wire \efuse_out[174] ;
 wire \efuse_out[175] ;
 wire \efuse_out[176] ;
 wire \efuse_out[177] ;
 wire \efuse_out[178] ;
 wire \efuse_out[179] ;
 wire \efuse_out[17] ;
 wire \efuse_out[180] ;
 wire \efuse_out[181] ;
 wire \efuse_out[182] ;
 wire \efuse_out[183] ;
 wire \efuse_out[184] ;
 wire \efuse_out[185] ;
 wire \efuse_out[186] ;
 wire \efuse_out[187] ;
 wire \efuse_out[188] ;
 wire \efuse_out[189] ;
 wire \efuse_out[18] ;
 wire \efuse_out[190] ;
 wire \efuse_out[191] ;
 wire \efuse_out[192] ;
 wire \efuse_out[193] ;
 wire \efuse_out[194] ;
 wire \efuse_out[195] ;
 wire \efuse_out[196] ;
 wire \efuse_out[197] ;
 wire \efuse_out[198] ;
 wire \efuse_out[199] ;
 wire \efuse_out[19] ;
 wire \efuse_out[1] ;
 wire \efuse_out[200] ;
 wire \efuse_out[201] ;
 wire \efuse_out[202] ;
 wire \efuse_out[203] ;
 wire \efuse_out[204] ;
 wire \efuse_out[205] ;
 wire \efuse_out[206] ;
 wire \efuse_out[207] ;
 wire \efuse_out[208] ;
 wire \efuse_out[209] ;
 wire \efuse_out[20] ;
 wire \efuse_out[210] ;
 wire \efuse_out[211] ;
 wire \efuse_out[212] ;
 wire \efuse_out[213] ;
 wire \efuse_out[214] ;
 wire \efuse_out[215] ;
 wire \efuse_out[216] ;
 wire \efuse_out[217] ;
 wire \efuse_out[218] ;
 wire \efuse_out[219] ;
 wire \efuse_out[21] ;
 wire \efuse_out[220] ;
 wire \efuse_out[221] ;
 wire \efuse_out[222] ;
 wire \efuse_out[223] ;
 wire \efuse_out[224] ;
 wire \efuse_out[225] ;
 wire \efuse_out[226] ;
 wire \efuse_out[227] ;
 wire \efuse_out[228] ;
 wire \efuse_out[229] ;
 wire \efuse_out[22] ;
 wire \efuse_out[230] ;
 wire \efuse_out[231] ;
 wire \efuse_out[232] ;
 wire \efuse_out[233] ;
 wire \efuse_out[234] ;
 wire \efuse_out[235] ;
 wire \efuse_out[236] ;
 wire \efuse_out[237] ;
 wire \efuse_out[238] ;
 wire \efuse_out[239] ;
 wire \efuse_out[23] ;
 wire \efuse_out[240] ;
 wire \efuse_out[241] ;
 wire \efuse_out[242] ;
 wire \efuse_out[243] ;
 wire \efuse_out[244] ;
 wire \efuse_out[245] ;
 wire \efuse_out[246] ;
 wire \efuse_out[247] ;
 wire \efuse_out[248] ;
 wire \efuse_out[249] ;
 wire \efuse_out[24] ;
 wire \efuse_out[250] ;
 wire \efuse_out[251] ;
 wire \efuse_out[252] ;
 wire \efuse_out[253] ;
 wire \efuse_out[254] ;
 wire \efuse_out[255] ;
 wire \efuse_out[256] ;
 wire \efuse_out[257] ;
 wire \efuse_out[258] ;
 wire \efuse_out[259] ;
 wire \efuse_out[25] ;
 wire \efuse_out[260] ;
 wire \efuse_out[261] ;
 wire \efuse_out[262] ;
 wire \efuse_out[263] ;
 wire \efuse_out[264] ;
 wire \efuse_out[265] ;
 wire \efuse_out[266] ;
 wire \efuse_out[267] ;
 wire \efuse_out[268] ;
 wire \efuse_out[269] ;
 wire \efuse_out[26] ;
 wire \efuse_out[270] ;
 wire \efuse_out[271] ;
 wire \efuse_out[272] ;
 wire \efuse_out[273] ;
 wire \efuse_out[274] ;
 wire \efuse_out[275] ;
 wire \efuse_out[276] ;
 wire \efuse_out[277] ;
 wire \efuse_out[278] ;
 wire \efuse_out[279] ;
 wire \efuse_out[27] ;
 wire \efuse_out[280] ;
 wire \efuse_out[281] ;
 wire \efuse_out[282] ;
 wire \efuse_out[283] ;
 wire \efuse_out[284] ;
 wire \efuse_out[285] ;
 wire \efuse_out[286] ;
 wire \efuse_out[287] ;
 wire \efuse_out[288] ;
 wire \efuse_out[289] ;
 wire \efuse_out[28] ;
 wire \efuse_out[290] ;
 wire \efuse_out[291] ;
 wire \efuse_out[292] ;
 wire \efuse_out[293] ;
 wire \efuse_out[294] ;
 wire \efuse_out[295] ;
 wire \efuse_out[296] ;
 wire \efuse_out[297] ;
 wire \efuse_out[298] ;
 wire \efuse_out[299] ;
 wire \efuse_out[29] ;
 wire \efuse_out[2] ;
 wire \efuse_out[300] ;
 wire \efuse_out[301] ;
 wire \efuse_out[302] ;
 wire \efuse_out[303] ;
 wire \efuse_out[304] ;
 wire \efuse_out[305] ;
 wire \efuse_out[306] ;
 wire \efuse_out[307] ;
 wire \efuse_out[308] ;
 wire \efuse_out[309] ;
 wire \efuse_out[30] ;
 wire \efuse_out[310] ;
 wire \efuse_out[311] ;
 wire \efuse_out[312] ;
 wire \efuse_out[313] ;
 wire \efuse_out[314] ;
 wire \efuse_out[315] ;
 wire \efuse_out[316] ;
 wire \efuse_out[317] ;
 wire \efuse_out[318] ;
 wire \efuse_out[319] ;
 wire \efuse_out[31] ;
 wire \efuse_out[320] ;
 wire \efuse_out[321] ;
 wire \efuse_out[322] ;
 wire \efuse_out[323] ;
 wire \efuse_out[324] ;
 wire \efuse_out[325] ;
 wire \efuse_out[326] ;
 wire \efuse_out[327] ;
 wire \efuse_out[328] ;
 wire \efuse_out[329] ;
 wire \efuse_out[32] ;
 wire \efuse_out[330] ;
 wire \efuse_out[331] ;
 wire \efuse_out[332] ;
 wire \efuse_out[333] ;
 wire \efuse_out[334] ;
 wire \efuse_out[335] ;
 wire \efuse_out[336] ;
 wire \efuse_out[337] ;
 wire \efuse_out[338] ;
 wire \efuse_out[339] ;
 wire \efuse_out[33] ;
 wire \efuse_out[340] ;
 wire \efuse_out[341] ;
 wire \efuse_out[342] ;
 wire \efuse_out[343] ;
 wire \efuse_out[344] ;
 wire \efuse_out[345] ;
 wire \efuse_out[346] ;
 wire \efuse_out[347] ;
 wire \efuse_out[348] ;
 wire \efuse_out[349] ;
 wire \efuse_out[34] ;
 wire \efuse_out[350] ;
 wire \efuse_out[351] ;
 wire \efuse_out[352] ;
 wire \efuse_out[353] ;
 wire \efuse_out[354] ;
 wire \efuse_out[355] ;
 wire \efuse_out[356] ;
 wire \efuse_out[357] ;
 wire \efuse_out[358] ;
 wire \efuse_out[359] ;
 wire \efuse_out[35] ;
 wire \efuse_out[360] ;
 wire \efuse_out[361] ;
 wire \efuse_out[362] ;
 wire \efuse_out[363] ;
 wire \efuse_out[364] ;
 wire \efuse_out[365] ;
 wire \efuse_out[366] ;
 wire \efuse_out[367] ;
 wire \efuse_out[368] ;
 wire \efuse_out[369] ;
 wire \efuse_out[36] ;
 wire \efuse_out[370] ;
 wire \efuse_out[371] ;
 wire \efuse_out[372] ;
 wire \efuse_out[373] ;
 wire \efuse_out[374] ;
 wire \efuse_out[375] ;
 wire \efuse_out[376] ;
 wire \efuse_out[377] ;
 wire \efuse_out[378] ;
 wire \efuse_out[379] ;
 wire \efuse_out[37] ;
 wire \efuse_out[380] ;
 wire \efuse_out[381] ;
 wire \efuse_out[382] ;
 wire \efuse_out[383] ;
 wire \efuse_out[384] ;
 wire \efuse_out[385] ;
 wire \efuse_out[386] ;
 wire \efuse_out[387] ;
 wire \efuse_out[388] ;
 wire \efuse_out[389] ;
 wire \efuse_out[38] ;
 wire \efuse_out[390] ;
 wire \efuse_out[391] ;
 wire \efuse_out[392] ;
 wire \efuse_out[393] ;
 wire \efuse_out[394] ;
 wire \efuse_out[395] ;
 wire \efuse_out[396] ;
 wire \efuse_out[397] ;
 wire \efuse_out[398] ;
 wire \efuse_out[399] ;
 wire \efuse_out[39] ;
 wire \efuse_out[3] ;
 wire \efuse_out[400] ;
 wire \efuse_out[401] ;
 wire \efuse_out[402] ;
 wire \efuse_out[403] ;
 wire \efuse_out[404] ;
 wire \efuse_out[405] ;
 wire \efuse_out[406] ;
 wire \efuse_out[407] ;
 wire \efuse_out[408] ;
 wire \efuse_out[409] ;
 wire \efuse_out[40] ;
 wire \efuse_out[410] ;
 wire \efuse_out[411] ;
 wire \efuse_out[412] ;
 wire \efuse_out[413] ;
 wire \efuse_out[414] ;
 wire \efuse_out[415] ;
 wire \efuse_out[416] ;
 wire \efuse_out[417] ;
 wire \efuse_out[418] ;
 wire \efuse_out[419] ;
 wire \efuse_out[41] ;
 wire \efuse_out[420] ;
 wire \efuse_out[421] ;
 wire \efuse_out[422] ;
 wire \efuse_out[423] ;
 wire \efuse_out[424] ;
 wire \efuse_out[425] ;
 wire \efuse_out[426] ;
 wire \efuse_out[427] ;
 wire \efuse_out[428] ;
 wire \efuse_out[429] ;
 wire \efuse_out[42] ;
 wire \efuse_out[430] ;
 wire \efuse_out[431] ;
 wire \efuse_out[432] ;
 wire \efuse_out[433] ;
 wire \efuse_out[434] ;
 wire \efuse_out[435] ;
 wire \efuse_out[436] ;
 wire \efuse_out[437] ;
 wire \efuse_out[438] ;
 wire \efuse_out[439] ;
 wire \efuse_out[43] ;
 wire \efuse_out[440] ;
 wire \efuse_out[441] ;
 wire \efuse_out[442] ;
 wire \efuse_out[443] ;
 wire \efuse_out[444] ;
 wire \efuse_out[445] ;
 wire \efuse_out[446] ;
 wire \efuse_out[447] ;
 wire \efuse_out[448] ;
 wire \efuse_out[449] ;
 wire \efuse_out[44] ;
 wire \efuse_out[450] ;
 wire \efuse_out[451] ;
 wire \efuse_out[452] ;
 wire \efuse_out[453] ;
 wire \efuse_out[454] ;
 wire \efuse_out[455] ;
 wire \efuse_out[456] ;
 wire \efuse_out[457] ;
 wire \efuse_out[458] ;
 wire \efuse_out[459] ;
 wire \efuse_out[45] ;
 wire \efuse_out[460] ;
 wire \efuse_out[461] ;
 wire \efuse_out[462] ;
 wire \efuse_out[463] ;
 wire \efuse_out[464] ;
 wire \efuse_out[465] ;
 wire \efuse_out[466] ;
 wire \efuse_out[467] ;
 wire \efuse_out[468] ;
 wire \efuse_out[469] ;
 wire \efuse_out[46] ;
 wire \efuse_out[470] ;
 wire \efuse_out[471] ;
 wire \efuse_out[472] ;
 wire \efuse_out[473] ;
 wire \efuse_out[474] ;
 wire \efuse_out[475] ;
 wire \efuse_out[476] ;
 wire \efuse_out[477] ;
 wire \efuse_out[478] ;
 wire \efuse_out[479] ;
 wire \efuse_out[47] ;
 wire \efuse_out[480] ;
 wire \efuse_out[481] ;
 wire \efuse_out[482] ;
 wire \efuse_out[483] ;
 wire \efuse_out[484] ;
 wire \efuse_out[485] ;
 wire \efuse_out[486] ;
 wire \efuse_out[487] ;
 wire \efuse_out[488] ;
 wire \efuse_out[489] ;
 wire \efuse_out[48] ;
 wire \efuse_out[490] ;
 wire \efuse_out[491] ;
 wire \efuse_out[492] ;
 wire \efuse_out[493] ;
 wire \efuse_out[494] ;
 wire \efuse_out[495] ;
 wire \efuse_out[496] ;
 wire \efuse_out[497] ;
 wire \efuse_out[498] ;
 wire \efuse_out[499] ;
 wire \efuse_out[49] ;
 wire \efuse_out[4] ;
 wire \efuse_out[500] ;
 wire \efuse_out[501] ;
 wire \efuse_out[502] ;
 wire \efuse_out[503] ;
 wire \efuse_out[504] ;
 wire \efuse_out[505] ;
 wire \efuse_out[506] ;
 wire \efuse_out[507] ;
 wire \efuse_out[508] ;
 wire \efuse_out[509] ;
 wire \efuse_out[50] ;
 wire \efuse_out[510] ;
 wire \efuse_out[511] ;
 wire \efuse_out[51] ;
 wire \efuse_out[52] ;
 wire \efuse_out[53] ;
 wire \efuse_out[54] ;
 wire \efuse_out[55] ;
 wire \efuse_out[56] ;
 wire \efuse_out[57] ;
 wire \efuse_out[58] ;
 wire \efuse_out[59] ;
 wire \efuse_out[5] ;
 wire \efuse_out[60] ;
 wire \efuse_out[61] ;
 wire \efuse_out[62] ;
 wire \efuse_out[63] ;
 wire \efuse_out[64] ;
 wire \efuse_out[65] ;
 wire \efuse_out[66] ;
 wire \efuse_out[67] ;
 wire \efuse_out[68] ;
 wire \efuse_out[69] ;
 wire \efuse_out[6] ;
 wire \efuse_out[70] ;
 wire \efuse_out[71] ;
 wire \efuse_out[72] ;
 wire \efuse_out[73] ;
 wire \efuse_out[74] ;
 wire \efuse_out[75] ;
 wire \efuse_out[76] ;
 wire \efuse_out[77] ;
 wire \efuse_out[78] ;
 wire \efuse_out[79] ;
 wire \efuse_out[7] ;
 wire \efuse_out[80] ;
 wire \efuse_out[81] ;
 wire \efuse_out[82] ;
 wire \efuse_out[83] ;
 wire \efuse_out[84] ;
 wire \efuse_out[85] ;
 wire \efuse_out[86] ;
 wire \efuse_out[87] ;
 wire \efuse_out[88] ;
 wire \efuse_out[89] ;
 wire \efuse_out[8] ;
 wire \efuse_out[90] ;
 wire \efuse_out[91] ;
 wire \efuse_out[92] ;
 wire \efuse_out[93] ;
 wire \efuse_out[94] ;
 wire \efuse_out[95] ;
 wire \efuse_out[96] ;
 wire \efuse_out[97] ;
 wire \efuse_out[98] ;
 wire \efuse_out[99] ;
 wire \efuse_out[9] ;
 wire one;
 wire \preset_n[0] ;
 wire \preset_n[10] ;
 wire \preset_n[11] ;
 wire \preset_n[12] ;
 wire \preset_n[13] ;
 wire \preset_n[14] ;
 wire \preset_n[15] ;
 wire \preset_n[1] ;
 wire \preset_n[2] ;
 wire \preset_n[3] ;
 wire \preset_n[4] ;
 wire \preset_n[5] ;
 wire \preset_n[6] ;
 wire \preset_n[7] ;
 wire \preset_n[8] ;
 wire \preset_n[9] ;
 wire \preset_n_reg[0] ;
 wire \preset_n_reg[10] ;
 wire \preset_n_reg[11] ;
 wire \preset_n_reg[12] ;
 wire \preset_n_reg[13] ;
 wire \preset_n_reg[14] ;
 wire \preset_n_reg[15] ;
 wire \preset_n_reg[1] ;
 wire \preset_n_reg[2] ;
 wire \preset_n_reg[3] ;
 wire \preset_n_reg[4] ;
 wire \preset_n_reg[5] ;
 wire \preset_n_reg[6] ;
 wire \preset_n_reg[7] ;
 wire \preset_n_reg[8] ;
 wire \preset_n_reg[9] ;
 wire \sense[0] ;
 wire \sense[10] ;
 wire \sense[11] ;
 wire \sense[12] ;
 wire \sense[13] ;
 wire \sense[14] ;
 wire \sense[15] ;
 wire \sense[1] ;
 wire \sense[2] ;
 wire \sense[3] ;
 wire \sense[4] ;
 wire \sense[5] ;
 wire \sense[6] ;
 wire \sense[7] ;
 wire \sense[8] ;
 wire \sense[9] ;
 wire \sense_del[0] ;
 wire \sense_del[10] ;
 wire \sense_del[11] ;
 wire \sense_del[12] ;
 wire \sense_del[13] ;
 wire \sense_del[14] ;
 wire \sense_del[15] ;
 wire \sense_del[1] ;
 wire \sense_del[2] ;
 wire \sense_del[3] ;
 wire \sense_del[4] ;
 wire \sense_del[5] ;
 wire \sense_del[6] ;
 wire \sense_del[7] ;
 wire \sense_del[8] ;
 wire \sense_del[9] ;
 wire \sense_reg[0] ;
 wire \sense_reg[10] ;
 wire \sense_reg[11] ;
 wire \sense_reg[12] ;
 wire \sense_reg[13] ;
 wire \sense_reg[14] ;
 wire \sense_reg[15] ;
 wire \sense_reg[1] ;
 wire \sense_reg[2] ;
 wire \sense_reg[3] ;
 wire \sense_reg[4] ;
 wire \sense_reg[5] ;
 wire \sense_reg[6] ;
 wire \sense_reg[7] ;
 wire \sense_reg[8] ;
 wire \sense_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2784_ (.I(net282),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2785_ (.I(\col_prog_n_reg[135] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2786_ (.I(\col_prog_n_reg[134] ),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(\col_prog_n_reg[133] ),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2788_ (.I(\col_prog_n_reg[132] ),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2789_ (.I(\col_prog_n_reg[131] ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2790_ (.I(\col_prog_n_reg[130] ),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2791_ (.I(\col_prog_n_reg[129] ),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2792_ (.I(\col_prog_n_reg[128] ),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2793_ (.I(\col_prog_n_reg[103] ),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2794_ (.I(\col_prog_n_reg[102] ),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2795_ (.I(\col_prog_n_reg[101] ),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2796_ (.I(\col_prog_n_reg[100] ),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2797_ (.I(\col_prog_n_reg[99] ),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2798_ (.I(\col_prog_n_reg[98] ),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2799_ (.I(\col_prog_n_reg[97] ),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2800_ (.I(\col_prog_n_reg[96] ),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2801_ (.I(\bit_sel_reg[46] ),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2802_ (.I(\bit_sel_reg[45] ),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2803_ (.I(\bit_sel_reg[14] ),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2804_ (.I(\bit_sel_reg[13] ),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2805_ (.I(\counter[8] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2806_ (.I(\counter[6] ),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2807_ (.I(\counter[5] ),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2808_ (.I(\counter[4] ),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2809_ (.I(\counter[3] ),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2810_ (.I(net285),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2811_ (.I(net66),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2812_ (.I(net65),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2813_ (.I(net64),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2814_ (.I(net62),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2815_ (.I(net61),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2816_ (.I(net58),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2817_ (.I(net57),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2818_ (.I(net56),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2819_ (.I(net54),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2820_ (.I(net83),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2821_ (.I(net78),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2822_ (.I(net52),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(\sense_reg[8] ),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2824_ (.I(\col_prog_n_reg[390] ),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2825_ (.I(\col_prog_n_reg[389] ),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(\col_prog_n_reg[388] ),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2827_ (.I(\col_prog_n_reg[387] ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2828_ (.I(\col_prog_n_reg[386] ),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2829_ (.I(\col_prog_n_reg[385] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2830_ (.I(\col_prog_n_reg[384] ),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2831_ (.I(\col_prog_n_reg[358] ),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2832_ (.I(\col_prog_n_reg[357] ),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2833_ (.I(\col_prog_n_reg[356] ),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2834_ (.I(\col_prog_n_reg[355] ),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2835_ (.I(\col_prog_n_reg[354] ),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2836_ (.I(\col_prog_n_reg[353] ),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2837_ (.I(\col_prog_n_reg[352] ),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2838_ (.I(\state[0] ),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2839_ (.I(net50),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _2840_ (.I(net361),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _2841_ (.I(net8),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _2842_ (.I(net355),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _2843_ (.I(net7),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2844_ (.I(net1),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2845_ (.I(net2),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2846_ (.I(net5),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2847_ (.I(net359),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2848_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2849_ (.A1(\counter[2] ),
    .A2(\counter[1] ),
    .A3(\counter[0] ),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2850_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .A4(\counter[0] ),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2851_ (.A1(_1334_),
    .A2(_1373_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(_1333_),
    .A2(_1374_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2853_ (.A1(\counter[5] ),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2854_ (.A1(_1332_),
    .A2(_1333_),
    .A3(_1374_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2855_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2856_ (.A1(_1332_),
    .A2(_1333_),
    .A3(_1374_),
    .A4(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2857_ (.A1(_1332_),
    .A2(_1333_),
    .A3(_1374_),
    .A4(_1379_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2858_ (.A1(\counter[9] ),
    .A2(\counter[8] ),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2859_ (.A1(_1380_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2860_ (.A1(\state[3] ),
    .A2(_1380_),
    .A3(_1382_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2861_ (.A1(\state[3] ),
    .A2(_1383_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2862_ (.A1(net7),
    .A2(net8),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2863_ (.A1(_1366_),
    .A2(_1368_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2864_ (.A1(net360),
    .A2(net347),
    .A3(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2865_ (.A1(net354),
    .A2(net9),
    .A3(net345),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2866_ (.A1(_1309_),
    .A2(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2867_ (.A1(\state[3] ),
    .A2(_1388_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2868_ (.A1(net48),
    .A2(net29),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2869_ (.A1(net186),
    .A2(net339),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2870_ (.A1(\col_prog_n_reg[153] ),
    .A2(net186),
    .B(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2871_ (.A1(net122),
    .A2(_1394_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2872_ (.A1(net48),
    .A2(net28),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2873_ (.A1(net186),
    .A2(net337),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2874_ (.A1(\col_prog_n_reg[152] ),
    .A2(net186),
    .B(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2875_ (.A1(net122),
    .A2(_1397_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2876_ (.A1(net47),
    .A2(net27),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2877_ (.A1(net186),
    .A2(net335),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2878_ (.A1(\col_prog_n_reg[151] ),
    .A2(net186),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2879_ (.A1(net122),
    .A2(_1400_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2880_ (.A1(net47),
    .A2(net26),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2881_ (.A1(net186),
    .A2(net333),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2882_ (.A1(\col_prog_n_reg[150] ),
    .A2(net186),
    .B(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2883_ (.A1(net122),
    .A2(_1403_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2884_ (.A1(net47),
    .A2(net25),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2885_ (.A1(net186),
    .A2(net331),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2886_ (.A1(\col_prog_n_reg[149] ),
    .A2(net186),
    .B(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2887_ (.A1(net122),
    .A2(_1406_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2888_ (.A1(net47),
    .A2(net24),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2889_ (.A1(net186),
    .A2(net330),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2890_ (.A1(\col_prog_n_reg[148] ),
    .A2(net186),
    .B(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2891_ (.A1(net122),
    .A2(_1409_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2892_ (.A1(net47),
    .A2(net22),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2893_ (.A1(net186),
    .A2(net327),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2894_ (.A1(\col_prog_n_reg[147] ),
    .A2(net186),
    .B(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2895_ (.A1(net122),
    .A2(_1412_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2896_ (.A1(net47),
    .A2(net21),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(net186),
    .A2(net325),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2898_ (.A1(\col_prog_n_reg[146] ),
    .A2(net186),
    .B(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2899_ (.A1(net122),
    .A2(_1415_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2900_ (.A1(net47),
    .A2(net20),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2901_ (.A1(net186),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2902_ (.A1(\col_prog_n_reg[145] ),
    .A2(net186),
    .B(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(net122),
    .A2(_1418_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2904_ (.A1(net47),
    .A2(net19),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2905_ (.A1(_1390_),
    .A2(net322),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2906_ (.A1(\col_prog_n_reg[144] ),
    .A2(_1390_),
    .B(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(_1385_),
    .A2(_1421_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2908_ (.A1(net46),
    .A2(net18),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2909_ (.A1(_1390_),
    .A2(net320),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2910_ (.A1(\col_prog_n_reg[143] ),
    .A2(_1390_),
    .B(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2911_ (.A1(_1385_),
    .A2(_1424_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2912_ (.A1(net46),
    .A2(net17),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2913_ (.A1(net187),
    .A2(net318),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2914_ (.A1(\col_prog_n_reg[142] ),
    .A2(net187),
    .B(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2915_ (.A1(net122),
    .A2(_1427_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2916_ (.A1(net46),
    .A2(net16),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2917_ (.A1(net187),
    .A2(net316),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2918_ (.A1(\col_prog_n_reg[141] ),
    .A2(net187),
    .B(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2919_ (.A1(net122),
    .A2(_1430_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2920_ (.A1(net46),
    .A2(net15),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2921_ (.A1(net187),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2922_ (.A1(\col_prog_n_reg[140] ),
    .A2(net187),
    .B(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2923_ (.A1(net122),
    .A2(_1433_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2924_ (.A1(net46),
    .A2(net14),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2925_ (.A1(net187),
    .A2(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2926_ (.A1(\col_prog_n_reg[139] ),
    .A2(net187),
    .B(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2927_ (.A1(net122),
    .A2(_1436_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2928_ (.A1(net46),
    .A2(net13),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2929_ (.A1(net187),
    .A2(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2930_ (.A1(\col_prog_n_reg[138] ),
    .A2(net187),
    .B(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2931_ (.A1(net122),
    .A2(_1439_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2932_ (.A1(net46),
    .A2(net43),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2933_ (.A1(net187),
    .A2(net308),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2934_ (.A1(\col_prog_n_reg[137] ),
    .A2(net187),
    .B(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2935_ (.A1(net122),
    .A2(_1442_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2936_ (.A1(net46),
    .A2(net42),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2937_ (.A1(net187),
    .A2(net305),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2938_ (.A1(\col_prog_n_reg[136] ),
    .A2(net187),
    .B(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(net122),
    .A2(_1445_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2940_ (.A1(_1384_),
    .A2(_1390_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2941_ (.A1(\counter[9] ),
    .A2(\counter[8] ),
    .A3(_1381_),
    .B(\state[3] ),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2942_ (.A1(net45),
    .A2(net41),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2943_ (.A1(net45),
    .A2(net41),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2944_ (.A1(net166),
    .A2(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2945_ (.A1(_1310_),
    .A2(_1446_),
    .B1(_1450_),
    .B2(net188),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2946_ (.A1(net45),
    .A2(net40),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2947_ (.A1(net45),
    .A2(net40),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2948_ (.A1(_1383_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2949_ (.A1(_1311_),
    .A2(_1446_),
    .B1(_1453_),
    .B2(_1390_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2950_ (.A1(net45),
    .A2(net39),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2951_ (.A1(net45),
    .A2(net39),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2952_ (.A1(_1383_),
    .A2(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2953_ (.A1(_1312_),
    .A2(_1446_),
    .B1(_1456_),
    .B2(_1390_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2954_ (.A1(net45),
    .A2(net38),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2955_ (.A1(net45),
    .A2(net38),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2956_ (.A1(_1383_),
    .A2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2957_ (.A1(_1313_),
    .A2(_1446_),
    .B1(net110),
    .B2(_1390_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2958_ (.A1(net45),
    .A2(net37),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2959_ (.A1(net45),
    .A2(net37),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2960_ (.A1(_1383_),
    .A2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2961_ (.A1(_1314_),
    .A2(_1446_),
    .B1(_1462_),
    .B2(_1390_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2962_ (.A1(net45),
    .A2(net34),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2963_ (.A1(net45),
    .A2(net34),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2964_ (.A1(net166),
    .A2(_1464_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2965_ (.A1(_1315_),
    .A2(_1446_),
    .B1(_1465_),
    .B2(net188),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2966_ (.A1(net45),
    .A2(net23),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2967_ (.A1(net45),
    .A2(net23),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2968_ (.A1(_1383_),
    .A2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2969_ (.A1(_1316_),
    .A2(_1446_),
    .B1(_1468_),
    .B2(_1390_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2970_ (.A1(net45),
    .A2(net12),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2971_ (.A1(net45),
    .A2(net12),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2972_ (.A1(_1383_),
    .A2(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2973_ (.A1(_1317_),
    .A2(_1446_),
    .B1(_1471_),
    .B2(_1390_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2974_ (.A1(net8),
    .A2(net7),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2975_ (.A1(net8),
    .A2(net7),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2976_ (.A1(net360),
    .A2(net9),
    .A3(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2977_ (.I(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2978_ (.A1(\state[3] ),
    .A2(_1474_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2979_ (.A1(\state[3] ),
    .A2(_1474_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2980_ (.A1(net48),
    .A2(net36),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2981_ (.A1(_1476_),
    .A2(net299),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2982_ (.A1(\col_prog_n_reg[127] ),
    .A2(_1476_),
    .B(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2983_ (.A1(net122),
    .A2(_1480_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2984_ (.A1(net48),
    .A2(net35),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2985_ (.A1(_1476_),
    .A2(net297),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2986_ (.A1(\col_prog_n_reg[126] ),
    .A2(_1476_),
    .B(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2987_ (.A1(net122),
    .A2(_1483_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2988_ (.A1(net48),
    .A2(net33),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2989_ (.A1(_1476_),
    .A2(net295),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2990_ (.A1(\col_prog_n_reg[125] ),
    .A2(_1476_),
    .B(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2991_ (.A1(net122),
    .A2(_1486_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2992_ (.A1(net48),
    .A2(net32),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2993_ (.A1(_1476_),
    .A2(net294),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2994_ (.A1(\col_prog_n_reg[124] ),
    .A2(_1476_),
    .B(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2995_ (.A1(net122),
    .A2(_1489_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2996_ (.A1(net48),
    .A2(net31),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2997_ (.A1(_1476_),
    .A2(net291),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2998_ (.A1(\col_prog_n_reg[123] ),
    .A2(_1476_),
    .B(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2999_ (.A1(net122),
    .A2(_1492_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3000_ (.A1(net48),
    .A2(net30),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3001_ (.A1(_1476_),
    .A2(net289),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3002_ (.A1(\col_prog_n_reg[122] ),
    .A2(_1476_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3003_ (.A1(net122),
    .A2(_1495_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3004_ (.A1(\col_prog_n_reg[121] ),
    .A2(net185),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3005_ (.A1(net339),
    .A2(net185),
    .B(_1496_),
    .C(net122),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3006_ (.A1(\col_prog_n_reg[120] ),
    .A2(net185),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3007_ (.A1(net337),
    .A2(net185),
    .B(_1497_),
    .C(net122),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3008_ (.A1(\col_prog_n_reg[119] ),
    .A2(net185),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3009_ (.A1(net335),
    .A2(net185),
    .B(_1498_),
    .C(net122),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3010_ (.A1(\col_prog_n_reg[118] ),
    .A2(net185),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3011_ (.A1(net333),
    .A2(net185),
    .B(_1499_),
    .C(net122),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3012_ (.A1(\col_prog_n_reg[117] ),
    .A2(net185),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3013_ (.A1(net331),
    .A2(net185),
    .B(_1500_),
    .C(net122),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3014_ (.A1(\col_prog_n_reg[116] ),
    .A2(net185),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3015_ (.A1(net330),
    .A2(net185),
    .B(_1501_),
    .C(net122),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3016_ (.A1(\col_prog_n_reg[115] ),
    .A2(net185),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3017_ (.A1(net327),
    .A2(net185),
    .B(_1502_),
    .C(net122),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3018_ (.A1(net325),
    .A2(_1476_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3019_ (.A1(\col_prog_n_reg[114] ),
    .A2(_1476_),
    .B(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3020_ (.A1(net122),
    .A2(_1504_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3021_ (.A1(_1416_),
    .A2(_1476_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3022_ (.A1(\col_prog_n_reg[113] ),
    .A2(_1476_),
    .B(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3023_ (.A1(net122),
    .A2(_1506_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3024_ (.A1(net322),
    .A2(_1476_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3025_ (.A1(\col_prog_n_reg[112] ),
    .A2(_1476_),
    .B(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3026_ (.A1(net122),
    .A2(_1508_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3027_ (.A1(\col_prog_n_reg[111] ),
    .A2(net185),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3028_ (.A1(net320),
    .A2(net185),
    .B(_1509_),
    .C(net122),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3029_ (.A1(\col_prog_n_reg[110] ),
    .A2(_1477_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3030_ (.A1(net318),
    .A2(_1477_),
    .B(_1510_),
    .C(net122),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3031_ (.A1(\col_prog_n_reg[109] ),
    .A2(_1477_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3032_ (.A1(net316),
    .A2(_1477_),
    .B(_1511_),
    .C(net122),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3033_ (.A1(\col_prog_n_reg[108] ),
    .A2(_1477_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3034_ (.A1(_1431_),
    .A2(_1477_),
    .B(_1512_),
    .C(net122),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3035_ (.A1(\col_prog_n_reg[107] ),
    .A2(_1477_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3036_ (.A1(_1434_),
    .A2(_1477_),
    .B(_1513_),
    .C(net122),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3037_ (.A1(\col_prog_n_reg[106] ),
    .A2(_1477_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3038_ (.A1(_1437_),
    .A2(_1477_),
    .B(_1514_),
    .C(net122),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3039_ (.A1(\col_prog_n_reg[105] ),
    .A2(_1477_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3040_ (.A1(net308),
    .A2(_1477_),
    .B(_1515_),
    .C(net122),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3041_ (.A1(\col_prog_n_reg[104] ),
    .A2(_1477_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3042_ (.A1(net305),
    .A2(_1477_),
    .B(_1516_),
    .C(net122),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3043_ (.A1(_1384_),
    .A2(_1476_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3044_ (.A1(net8),
    .A2(net9),
    .A3(net7),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3045_ (.A1(net354),
    .A2(net286),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3046_ (.A1(net354),
    .A2(net286),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3047_ (.A1(_1449_),
    .A2(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3048_ (.A1(_1383_),
    .A2(_1477_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3049_ (.A1(_1318_),
    .A2(_1517_),
    .B1(_1521_),
    .B2(_1522_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3050_ (.A1(_1452_),
    .A2(_1520_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3051_ (.A1(_1319_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1523_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3052_ (.A1(_1455_),
    .A2(_1520_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3053_ (.A1(_1320_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1524_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3054_ (.A1(_1458_),
    .A2(_1520_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3055_ (.A1(_1321_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1525_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3056_ (.A1(_1461_),
    .A2(_1520_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3057_ (.A1(_1322_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1526_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3058_ (.A1(_1464_),
    .A2(_1520_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3059_ (.A1(_1323_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1527_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3060_ (.A1(_1467_),
    .A2(_1520_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3061_ (.A1(_1324_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1528_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3062_ (.A1(_1470_),
    .A2(_1520_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3063_ (.A1(_1325_),
    .A2(_1517_),
    .B1(_1522_),
    .B2(_1529_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3064_ (.A1(net7),
    .A2(_1366_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3065_ (.A1(net8),
    .A2(net348),
    .A3(_1368_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3066_ (.A1(net360),
    .A2(net271),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3067_ (.A1(net353),
    .A2(net8),
    .A3(net348),
    .A4(_1368_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3068_ (.A1(_1309_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3069_ (.A1(\state[3] ),
    .A2(_1532_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3070_ (.A1(\col_prog_n_reg[95] ),
    .A2(net162),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3071_ (.A1(net299),
    .A2(net162),
    .B(_1536_),
    .C(net117),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3072_ (.A1(\col_prog_n_reg[94] ),
    .A2(net162),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3073_ (.A1(net297),
    .A2(net162),
    .B(_1537_),
    .C(net117),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3074_ (.A1(\col_prog_n_reg[93] ),
    .A2(net162),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3075_ (.A1(net295),
    .A2(net162),
    .B(_1538_),
    .C(net117),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3076_ (.A1(net294),
    .A2(net184),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3077_ (.A1(\col_prog_n_reg[92] ),
    .A2(net184),
    .B(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3078_ (.A1(net117),
    .A2(_1540_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3079_ (.A1(\col_prog_n_reg[91] ),
    .A2(net162),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3080_ (.A1(net291),
    .A2(net162),
    .B(_1541_),
    .C(net117),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3081_ (.A1(net289),
    .A2(net184),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3082_ (.A1(\col_prog_n_reg[90] ),
    .A2(net184),
    .B(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3083_ (.A1(net117),
    .A2(_1543_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3084_ (.A1(\col_prog_n_reg[89] ),
    .A2(net162),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3085_ (.A1(net339),
    .A2(net162),
    .B(_1544_),
    .C(net117),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3086_ (.A1(\col_prog_n_reg[88] ),
    .A2(net162),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3087_ (.A1(net337),
    .A2(net162),
    .B(_1545_),
    .C(net117),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3088_ (.A1(\col_prog_n_reg[87] ),
    .A2(net162),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3089_ (.A1(net335),
    .A2(net162),
    .B(_1546_),
    .C(net117),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3090_ (.A1(\col_prog_n_reg[86] ),
    .A2(net162),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3091_ (.A1(net333),
    .A2(net162),
    .B(_1547_),
    .C(net117),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3092_ (.A1(\col_prog_n_reg[85] ),
    .A2(net162),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3093_ (.A1(net331),
    .A2(net162),
    .B(_1548_),
    .C(net117),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3094_ (.A1(\col_prog_n_reg[84] ),
    .A2(net163),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3095_ (.A1(net330),
    .A2(net162),
    .B(_1549_),
    .C(net117),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3096_ (.A1(\col_prog_n_reg[83] ),
    .A2(net163),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3097_ (.A1(net327),
    .A2(net163),
    .B(_1550_),
    .C(net117),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3098_ (.A1(\col_prog_n_reg[82] ),
    .A2(net163),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3099_ (.A1(net325),
    .A2(net163),
    .B(_1551_),
    .C(net117),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3100_ (.A1(\col_prog_n_reg[81] ),
    .A2(net163),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3101_ (.A1(_1416_),
    .A2(net163),
    .B(_1552_),
    .C(net117),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3102_ (.A1(\col_prog_n_reg[80] ),
    .A2(net163),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3103_ (.A1(net322),
    .A2(net163),
    .B(_1553_),
    .C(net117),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3104_ (.A1(\col_prog_n_reg[79] ),
    .A2(net163),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3105_ (.A1(net320),
    .A2(net163),
    .B(_1554_),
    .C(net117),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3106_ (.A1(\col_prog_n_reg[78] ),
    .A2(net163),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3107_ (.A1(net318),
    .A2(net163),
    .B(_1555_),
    .C(net117),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3108_ (.A1(\col_prog_n_reg[77] ),
    .A2(net163),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3109_ (.A1(net316),
    .A2(net163),
    .B(_1556_),
    .C(net117),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3110_ (.A1(\col_prog_n_reg[76] ),
    .A2(_1535_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3111_ (.A1(_1431_),
    .A2(_1535_),
    .B(_1557_),
    .C(net117),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3112_ (.A1(\col_prog_n_reg[75] ),
    .A2(_1535_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3113_ (.A1(_1434_),
    .A2(_1535_),
    .B(_1558_),
    .C(net117),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3114_ (.A1(\col_prog_n_reg[74] ),
    .A2(_1535_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3115_ (.A1(_1437_),
    .A2(_1535_),
    .B(_1559_),
    .C(net117),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3116_ (.A1(\col_prog_n_reg[73] ),
    .A2(_1535_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3117_ (.A1(net308),
    .A2(_1535_),
    .B(_1560_),
    .C(net117),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3118_ (.A1(\col_prog_n_reg[72] ),
    .A2(_1535_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3119_ (.A1(net305),
    .A2(_1535_),
    .B(_1561_),
    .C(net117),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3120_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[71] ),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3121_ (.A1(_1521_),
    .A2(net270),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3122_ (.A1(net360),
    .A2(net288),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3123_ (.A1(net353),
    .A2(net287),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3124_ (.A1(net360),
    .A2(net288),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3125_ (.A1(\col_prog_n_reg[71] ),
    .A2(net269),
    .B1(_1563_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3126_ (.A1(_1562_),
    .A2(_1567_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3127_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[70] ),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3128_ (.A1(_1523_),
    .A2(net270),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3129_ (.A1(\col_prog_n_reg[70] ),
    .A2(net269),
    .B1(_1565_),
    .B2(_1569_),
    .C(net166),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3130_ (.A1(_1568_),
    .A2(_1570_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3131_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[69] ),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3132_ (.A1(_1524_),
    .A2(net270),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3133_ (.A1(\col_prog_n_reg[69] ),
    .A2(net269),
    .B1(_1565_),
    .B2(_1572_),
    .C(net166),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3134_ (.A1(_1571_),
    .A2(_1573_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3135_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[68] ),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3136_ (.A1(_1525_),
    .A2(net270),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3137_ (.A1(\col_prog_n_reg[68] ),
    .A2(net269),
    .B1(_1565_),
    .B2(_1575_),
    .C(net166),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3138_ (.A1(_1574_),
    .A2(_1576_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3139_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[67] ),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3140_ (.A1(_1526_),
    .A2(net270),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3141_ (.A1(\col_prog_n_reg[67] ),
    .A2(net269),
    .B1(_1565_),
    .B2(_1578_),
    .C(net166),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3142_ (.A1(_1577_),
    .A2(_1579_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3143_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[66] ),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3144_ (.A1(_1527_),
    .A2(net270),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3145_ (.A1(\col_prog_n_reg[66] ),
    .A2(net269),
    .B1(_1565_),
    .B2(_1581_),
    .C(net166),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3146_ (.A1(_1580_),
    .A2(_1582_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3147_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[65] ),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3148_ (.A1(_1528_),
    .A2(net270),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3149_ (.A1(\col_prog_n_reg[65] ),
    .A2(net269),
    .B1(net268),
    .B2(_1584_),
    .C(net166),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3150_ (.A1(_1583_),
    .A2(_1585_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3151_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[64] ),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3152_ (.A1(_1529_),
    .A2(net270),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3153_ (.A1(\col_prog_n_reg[64] ),
    .A2(net269),
    .B1(net268),
    .B2(_1587_),
    .C(net166),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3154_ (.A1(_1586_),
    .A2(_1588_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3155_ (.A1(_1368_),
    .A2(net8),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3156_ (.A1(_1366_),
    .A2(_1367_),
    .A3(net7),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3157_ (.A1(net360),
    .A2(net260),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3158_ (.A1(net354),
    .A2(net347),
    .A3(net262),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3159_ (.A1(\state[3] ),
    .A2(_1591_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3160_ (.A1(\col_prog_n_reg[63] ),
    .A2(net160),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3161_ (.A1(net299),
    .A2(net160),
    .B(_1594_),
    .C(net117),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3162_ (.A1(\col_prog_n_reg[62] ),
    .A2(net160),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3163_ (.A1(net297),
    .A2(net160),
    .B(_1595_),
    .C(net117),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3164_ (.A1(\col_prog_n_reg[61] ),
    .A2(net160),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3165_ (.A1(net295),
    .A2(net160),
    .B(_1596_),
    .C(net117),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3166_ (.A1(\col_prog_n_reg[60] ),
    .A2(net160),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3167_ (.A1(net294),
    .A2(net160),
    .B(_1597_),
    .C(net117),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3168_ (.A1(\col_prog_n_reg[59] ),
    .A2(net160),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3169_ (.A1(net291),
    .A2(net160),
    .B(_1598_),
    .C(net117),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3170_ (.A1(\col_prog_n_reg[58] ),
    .A2(net160),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3171_ (.A1(net289),
    .A2(net160),
    .B(_1599_),
    .C(net117),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3172_ (.A1(\col_prog_n_reg[57] ),
    .A2(net160),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3173_ (.A1(net339),
    .A2(net160),
    .B(_1600_),
    .C(net117),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3174_ (.A1(\col_prog_n_reg[56] ),
    .A2(net160),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3175_ (.A1(net337),
    .A2(net160),
    .B(_1601_),
    .C(net117),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3176_ (.A1(\col_prog_n_reg[55] ),
    .A2(net160),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3177_ (.A1(net335),
    .A2(net160),
    .B(_1602_),
    .C(net117),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3178_ (.A1(\col_prog_n_reg[54] ),
    .A2(net160),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3179_ (.A1(net333),
    .A2(net160),
    .B(_1603_),
    .C(net117),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3180_ (.A1(\col_prog_n_reg[53] ),
    .A2(net161),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3181_ (.A1(net331),
    .A2(net161),
    .B(_1604_),
    .C(net117),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3182_ (.A1(\col_prog_n_reg[52] ),
    .A2(net161),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3183_ (.A1(net330),
    .A2(net161),
    .B(_1605_),
    .C(net117),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3184_ (.A1(\col_prog_n_reg[51] ),
    .A2(net161),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3185_ (.A1(net327),
    .A2(net161),
    .B(_1606_),
    .C(net117),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3186_ (.A1(\col_prog_n_reg[50] ),
    .A2(net161),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3187_ (.A1(net325),
    .A2(net161),
    .B(_1607_),
    .C(net117),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3188_ (.A1(\col_prog_n_reg[49] ),
    .A2(net161),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3189_ (.A1(_1416_),
    .A2(net161),
    .B(_1608_),
    .C(net117),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3190_ (.A1(\col_prog_n_reg[48] ),
    .A2(net161),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3191_ (.A1(net322),
    .A2(net161),
    .B(_1609_),
    .C(net117),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3192_ (.A1(\col_prog_n_reg[47] ),
    .A2(net161),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3193_ (.A1(net320),
    .A2(net161),
    .B(_1610_),
    .C(net117),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3194_ (.A1(\col_prog_n_reg[46] ),
    .A2(net161),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3195_ (.A1(net318),
    .A2(net161),
    .B(_1611_),
    .C(net117),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3196_ (.A1(\col_prog_n_reg[45] ),
    .A2(_1593_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3197_ (.A1(net316),
    .A2(net161),
    .B(_1612_),
    .C(net117),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3198_ (.A1(\col_prog_n_reg[44] ),
    .A2(_1593_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3199_ (.A1(_1431_),
    .A2(_1593_),
    .B(_1613_),
    .C(net117),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3200_ (.A1(\col_prog_n_reg[43] ),
    .A2(_1593_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3201_ (.A1(_1434_),
    .A2(_1593_),
    .B(_1614_),
    .C(net117),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3202_ (.A1(\col_prog_n_reg[42] ),
    .A2(_1593_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3203_ (.A1(_1437_),
    .A2(_1593_),
    .B(_1615_),
    .C(net117),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3204_ (.A1(\col_prog_n_reg[41] ),
    .A2(_1593_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3205_ (.A1(net308),
    .A2(_1593_),
    .B(_1616_),
    .C(net117),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3206_ (.A1(\col_prog_n_reg[40] ),
    .A2(_1593_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3207_ (.A1(net305),
    .A2(_1593_),
    .B(_1617_),
    .C(net117),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3208_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[39] ),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3209_ (.A1(_1521_),
    .A2(net260),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3210_ (.A1(\col_prog_n_reg[39] ),
    .A2(_1592_),
    .B1(_1619_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3211_ (.A1(_1618_),
    .A2(_1620_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3212_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[38] ),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3213_ (.A1(_1523_),
    .A2(net260),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3214_ (.A1(\col_prog_n_reg[38] ),
    .A2(_1592_),
    .B1(_1622_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3215_ (.A1(_1621_),
    .A2(_1623_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3216_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[37] ),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3217_ (.A1(_1524_),
    .A2(net260),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3218_ (.A1(\col_prog_n_reg[37] ),
    .A2(_1592_),
    .B1(_1625_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3219_ (.A1(_1624_),
    .A2(_1626_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3220_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[36] ),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3221_ (.A1(_1525_),
    .A2(net260),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3222_ (.A1(\col_prog_n_reg[36] ),
    .A2(_1592_),
    .B1(_1628_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3223_ (.A1(_1627_),
    .A2(_1629_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3224_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[35] ),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3225_ (.A1(_1526_),
    .A2(net260),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3226_ (.A1(\col_prog_n_reg[35] ),
    .A2(_1592_),
    .B1(_1631_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3227_ (.A1(_1630_),
    .A2(_1632_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3228_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[34] ),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3229_ (.A1(_1527_),
    .A2(net260),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3230_ (.A1(\col_prog_n_reg[34] ),
    .A2(_1592_),
    .B1(_1634_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3231_ (.A1(_1633_),
    .A2(_1635_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3232_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[33] ),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3233_ (.A1(_1528_),
    .A2(net260),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3234_ (.A1(\col_prog_n_reg[33] ),
    .A2(_1592_),
    .B1(_1637_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3235_ (.A1(_1636_),
    .A2(_1638_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3236_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[32] ),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3237_ (.A1(_1529_),
    .A2(net260),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3238_ (.A1(\col_prog_n_reg[32] ),
    .A2(_1592_),
    .B1(_1640_),
    .B2(_1565_),
    .C(net166),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3239_ (.A1(_1639_),
    .A2(_1641_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3240_ (.A1(\state[3] ),
    .A2(_1519_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3241_ (.A1(\col_prog_n_reg[31] ),
    .A2(net182),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3242_ (.A1(net299),
    .A2(net182),
    .B(_1643_),
    .C(net117),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3243_ (.A1(\col_prog_n_reg[30] ),
    .A2(net182),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3244_ (.A1(net297),
    .A2(net182),
    .B(_1644_),
    .C(net117),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3245_ (.A1(\col_prog_n_reg[29] ),
    .A2(net182),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3246_ (.A1(net295),
    .A2(net182),
    .B(_1645_),
    .C(net117),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3247_ (.A1(\col_prog_n_reg[28] ),
    .A2(net182),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3248_ (.A1(net294),
    .A2(net182),
    .B(_1646_),
    .C(net117),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3249_ (.A1(\col_prog_n_reg[27] ),
    .A2(net182),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3250_ (.A1(net291),
    .A2(net182),
    .B(_1647_),
    .C(net117),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3251_ (.A1(\col_prog_n_reg[26] ),
    .A2(net182),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3252_ (.A1(net289),
    .A2(net182),
    .B(_1648_),
    .C(net117),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3253_ (.A1(\col_prog_n_reg[25] ),
    .A2(net182),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3254_ (.A1(net339),
    .A2(net182),
    .B(_1649_),
    .C(net117),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3255_ (.A1(\col_prog_n_reg[24] ),
    .A2(net182),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3256_ (.A1(net337),
    .A2(net182),
    .B(_1650_),
    .C(net117),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3257_ (.A1(\col_prog_n_reg[23] ),
    .A2(net182),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3258_ (.A1(net335),
    .A2(net182),
    .B(_1651_),
    .C(net117),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3259_ (.A1(\col_prog_n_reg[22] ),
    .A2(net182),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3260_ (.A1(net333),
    .A2(net182),
    .B(_1652_),
    .C(net117),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3261_ (.A1(\col_prog_n_reg[21] ),
    .A2(net182),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3262_ (.A1(net331),
    .A2(net182),
    .B(_1653_),
    .C(net117),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3263_ (.A1(\col_prog_n_reg[20] ),
    .A2(net182),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3264_ (.A1(net330),
    .A2(net182),
    .B(_1654_),
    .C(net117),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3265_ (.A1(\col_prog_n_reg[19] ),
    .A2(net182),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3266_ (.A1(net327),
    .A2(net182),
    .B(_1655_),
    .C(net117),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3267_ (.A1(\col_prog_n_reg[18] ),
    .A2(net182),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3268_ (.A1(net325),
    .A2(net182),
    .B(_1656_),
    .C(net117),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3269_ (.A1(\col_prog_n_reg[17] ),
    .A2(net183),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3270_ (.A1(_1416_),
    .A2(net183),
    .B(_1657_),
    .C(net117),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3271_ (.A1(\col_prog_n_reg[16] ),
    .A2(net183),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3272_ (.A1(net322),
    .A2(net183),
    .B(_1658_),
    .C(net117),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3273_ (.A1(\col_prog_n_reg[15] ),
    .A2(net183),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3274_ (.A1(net320),
    .A2(net183),
    .B(_1659_),
    .C(net117),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3275_ (.A1(\col_prog_n_reg[14] ),
    .A2(net183),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3276_ (.A1(net318),
    .A2(net183),
    .B(_1660_),
    .C(net117),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3277_ (.A1(\col_prog_n_reg[13] ),
    .A2(net183),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3278_ (.A1(net316),
    .A2(net183),
    .B(_1661_),
    .C(net117),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3279_ (.A1(\col_prog_n_reg[12] ),
    .A2(net183),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3280_ (.A1(_1431_),
    .A2(net183),
    .B(_1662_),
    .C(net117),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3281_ (.A1(\col_prog_n_reg[11] ),
    .A2(net183),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3282_ (.A1(_1434_),
    .A2(net183),
    .B(_1663_),
    .C(net117),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3283_ (.A1(\col_prog_n_reg[10] ),
    .A2(net183),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3284_ (.A1(_1437_),
    .A2(net183),
    .B(_1664_),
    .C(net117),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3285_ (.A1(\col_prog_n_reg[9] ),
    .A2(net183),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3286_ (.A1(net308),
    .A2(net183),
    .B(_1665_),
    .C(net117),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3287_ (.A1(\col_prog_n_reg[8] ),
    .A2(net183),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3288_ (.A1(net305),
    .A2(net183),
    .B(_1666_),
    .C(net117),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3289_ (.A1(\col_prog_n_reg[7] ),
    .A2(_1642_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3290_ (.A1(_1448_),
    .A2(_1642_),
    .B(_1667_),
    .C(net122),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3291_ (.A1(\col_prog_n_reg[6] ),
    .A2(_1642_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3292_ (.A1(_1451_),
    .A2(_1642_),
    .B(_1668_),
    .C(net122),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3293_ (.A1(\col_prog_n_reg[5] ),
    .A2(_1642_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3294_ (.A1(_1454_),
    .A2(_1642_),
    .B(_1669_),
    .C(net122),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3295_ (.A1(\col_prog_n_reg[4] ),
    .A2(_1642_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3296_ (.A1(_1457_),
    .A2(_1642_),
    .B(_1670_),
    .C(net122),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3297_ (.A1(\col_prog_n_reg[3] ),
    .A2(_1642_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3298_ (.A1(_1460_),
    .A2(_1642_),
    .B(_1671_),
    .C(net122),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3299_ (.A1(\col_prog_n_reg[2] ),
    .A2(_1642_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3300_ (.A1(_1463_),
    .A2(_1642_),
    .B(_1672_),
    .C(net122),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3301_ (.A1(\col_prog_n_reg[1] ),
    .A2(_1642_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3302_ (.A1(_1466_),
    .A2(_1642_),
    .B(_1673_),
    .C(net122),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3303_ (.A1(\col_prog_n_reg[0] ),
    .A2(net183),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3304_ (.A1(_1469_),
    .A2(net183),
    .B(_1674_),
    .C(net117),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3305_ (.A1(\state[0] ),
    .A2(\state[2] ),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3306_ (.A1(\state[0] ),
    .A2(\state[2] ),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3307_ (.A1(\bit_sel_reg[63] ),
    .A2(_1675_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3308_ (.A1(net1),
    .A2(net2),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3309_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3310_ (.I(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3311_ (.A1(net4),
    .A2(net5),
    .A3(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3312_ (.A1(net11),
    .A2(net49),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3313_ (.A1(net51),
    .A2(_1682_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3314_ (.A1(net50),
    .A2(_1683_),
    .B(\state[2] ),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3315_ (.I(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3316_ (.A1(net6),
    .A2(_1676_),
    .A3(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3317_ (.A1(_1681_),
    .A2(net100),
    .B(_1677_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(\bit_sel_reg[62] ),
    .A2(net259),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3319_ (.A1(net1),
    .A2(_1370_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3320_ (.A1(_1369_),
    .A2(net2),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3321_ (.A1(net3),
    .A2(_1688_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3322_ (.A1(net3),
    .A2(net4),
    .A3(_1688_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3323_ (.A1(_1371_),
    .A2(_1691_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3324_ (.A1(net100),
    .A2(_1692_),
    .B(_1687_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3325_ (.A1(\bit_sel_reg[61] ),
    .A2(_1675_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3326_ (.A1(_1369_),
    .A2(net2),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3327_ (.A1(net1),
    .A2(_1370_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3328_ (.A1(net3),
    .A2(_1694_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3329_ (.A1(net3),
    .A2(net4),
    .A3(_1694_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3330_ (.A1(_1371_),
    .A2(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3331_ (.A1(_1686_),
    .A2(_1698_),
    .B(_1693_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3332_ (.A1(\bit_sel_reg[60] ),
    .A2(net259),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3333_ (.A1(net1),
    .A2(net2),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3334_ (.A1(net3),
    .A2(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3335_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(_1700_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3336_ (.A1(_1686_),
    .A2(_1702_),
    .B(_1699_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(\bit_sel_reg[59] ),
    .A2(net258),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3338_ (.A1(net3),
    .A2(_1678_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3339_ (.A1(net4),
    .A2(net5),
    .A3(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3340_ (.A1(net99),
    .A2(_1705_),
    .B(_1703_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3341_ (.A1(\bit_sel_reg[58] ),
    .A2(net259),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3342_ (.A1(net3),
    .A2(_1689_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3343_ (.A1(net4),
    .A2(net5),
    .A3(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3344_ (.A1(_1686_),
    .A2(_1708_),
    .B(_1706_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3345_ (.A1(\bit_sel_reg[57] ),
    .A2(net259),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3346_ (.A1(net3),
    .A2(_1695_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3347_ (.A1(net4),
    .A2(net5),
    .A3(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3348_ (.A1(net100),
    .A2(_1711_),
    .B(_1709_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3349_ (.A1(\bit_sel_reg[56] ),
    .A2(net259),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3350_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3351_ (.A1(net4),
    .A2(net5),
    .A3(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3352_ (.A1(_1686_),
    .A2(_1714_),
    .B(_1712_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3353_ (.A1(\bit_sel_reg[55] ),
    .A2(_1675_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3354_ (.A1(net4),
    .A2(_1679_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3355_ (.A1(net5),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3356_ (.A1(net100),
    .A2(_1717_),
    .B(_1715_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3357_ (.A1(\bit_sel_reg[54] ),
    .A2(_1675_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3358_ (.A1(net4),
    .A2(_1690_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3359_ (.A1(net5),
    .A2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3360_ (.A1(_1686_),
    .A2(_1720_),
    .B(_1718_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3361_ (.A1(\bit_sel_reg[53] ),
    .A2(_1675_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3362_ (.A1(net4),
    .A2(_1696_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3363_ (.A1(net5),
    .A2(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3364_ (.A1(_1686_),
    .A2(_1723_),
    .B(_1721_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3365_ (.A1(\bit_sel_reg[52] ),
    .A2(_1675_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3366_ (.A1(net4),
    .A2(_1701_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3367_ (.A1(net5),
    .A2(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3368_ (.A1(net100),
    .A2(_1726_),
    .B(_1724_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3369_ (.A1(\bit_sel_reg[51] ),
    .A2(net258),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3370_ (.A1(net3),
    .A2(net4),
    .A3(_1678_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3371_ (.A1(net5),
    .A2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3372_ (.A1(net99),
    .A2(_1729_),
    .B(_1727_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3373_ (.A1(\bit_sel_reg[50] ),
    .A2(net258),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3374_ (.A1(net3),
    .A2(net4),
    .A3(_1689_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3375_ (.A1(net5),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3376_ (.A1(net99),
    .A2(_1732_),
    .B(_1730_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3377_ (.A1(\bit_sel_reg[49] ),
    .A2(_1675_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3378_ (.A1(net3),
    .A2(net4),
    .A3(_1695_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3379_ (.A1(net5),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3380_ (.A1(net100),
    .A2(_1735_),
    .B(_1733_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3381_ (.A1(\bit_sel_reg[48] ),
    .A2(net258),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3382_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .A4(net4),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3383_ (.A1(net5),
    .A2(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3384_ (.A1(net99),
    .A2(_1738_),
    .B(_1736_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3385_ (.A1(\bit_sel_reg[47] ),
    .A2(net259),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3386_ (.A1(net4),
    .A2(_1371_),
    .A3(_1680_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3387_ (.A1(net100),
    .A2(_1740_),
    .B(_1739_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3388_ (.A1(net5),
    .A2(net100),
    .A3(_1691_),
    .B1(_1676_),
    .B2(_1326_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3389_ (.A1(net5),
    .A2(_1686_),
    .A3(_1697_),
    .B1(_1676_),
    .B2(_1327_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3390_ (.A1(\bit_sel_reg[44] ),
    .A2(net259),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3391_ (.A1(net3),
    .A2(net4),
    .A3(_1371_),
    .A4(_1700_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3392_ (.A1(_1686_),
    .A2(_1742_),
    .B(_1741_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3393_ (.A1(\bit_sel_reg[43] ),
    .A2(net258),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3394_ (.A1(net4),
    .A2(_1371_),
    .A3(_1704_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3395_ (.A1(net99),
    .A2(_1744_),
    .B(_1743_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3396_ (.A1(\bit_sel_reg[42] ),
    .A2(net259),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3397_ (.A1(net4),
    .A2(_1371_),
    .A3(_1707_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3398_ (.A1(net100),
    .A2(_1746_),
    .B(_1745_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3399_ (.A1(\bit_sel_reg[41] ),
    .A2(net259),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3400_ (.A1(net4),
    .A2(_1371_),
    .A3(_1710_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3401_ (.A1(net100),
    .A2(_1748_),
    .B(_1747_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3402_ (.A1(\bit_sel_reg[40] ),
    .A2(net259),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3403_ (.A1(net4),
    .A2(_1371_),
    .A3(_1713_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3404_ (.A1(_1686_),
    .A2(_1750_),
    .B(_1749_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3405_ (.A1(\bit_sel_reg[39] ),
    .A2(_1675_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3406_ (.A1(_1371_),
    .A2(_1716_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3407_ (.A1(net100),
    .A2(_1752_),
    .B(_1751_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3408_ (.A1(\bit_sel_reg[38] ),
    .A2(_1675_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3409_ (.A1(_1371_),
    .A2(_1719_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3410_ (.A1(_1686_),
    .A2(_1754_),
    .B(_1753_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3411_ (.A1(\bit_sel_reg[37] ),
    .A2(_1675_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3412_ (.A1(_1371_),
    .A2(_1722_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3413_ (.A1(_1686_),
    .A2(_1756_),
    .B(_1755_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3414_ (.A1(\bit_sel_reg[36] ),
    .A2(_1675_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(_1371_),
    .A2(_1725_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3416_ (.A1(net100),
    .A2(_1758_),
    .B(_1757_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3417_ (.A1(\bit_sel_reg[35] ),
    .A2(net258),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3418_ (.A1(_1371_),
    .A2(_1728_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3419_ (.A1(net99),
    .A2(_1760_),
    .B(_1759_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3420_ (.A1(\bit_sel_reg[34] ),
    .A2(net258),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(_1371_),
    .A2(_1731_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3422_ (.A1(net99),
    .A2(_1762_),
    .B(_1761_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3423_ (.A1(\bit_sel_reg[33] ),
    .A2(_1675_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3424_ (.A1(_1371_),
    .A2(_1734_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3425_ (.A1(net100),
    .A2(_1764_),
    .B(_1763_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3426_ (.A1(\bit_sel_reg[32] ),
    .A2(net258),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3427_ (.A1(_1371_),
    .A2(_1737_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3428_ (.A1(net99),
    .A2(_1766_),
    .B(_1765_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3429_ (.A1(\bit_sel_reg[31] ),
    .A2(_1675_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3430_ (.A1(net6),
    .A2(_1675_),
    .A3(_1684_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3431_ (.A1(_1681_),
    .A2(net159),
    .B(_1767_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3432_ (.A1(\bit_sel_reg[30] ),
    .A2(net259),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3433_ (.A1(_1692_),
    .A2(net159),
    .B(_1769_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3434_ (.A1(\bit_sel_reg[29] ),
    .A2(_1675_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3435_ (.A1(_1698_),
    .A2(_1768_),
    .B(_1770_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3436_ (.A1(\bit_sel_reg[28] ),
    .A2(net259),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3437_ (.A1(_1702_),
    .A2(_1768_),
    .B(_1771_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(\bit_sel_reg[27] ),
    .A2(net258),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3439_ (.A1(_1705_),
    .A2(net159),
    .B(_1772_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3440_ (.A1(\bit_sel_reg[26] ),
    .A2(net259),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3441_ (.A1(_1708_),
    .A2(_1768_),
    .B(_1773_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3442_ (.A1(\bit_sel_reg[25] ),
    .A2(net259),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3443_ (.A1(_1711_),
    .A2(net159),
    .B(_1774_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3444_ (.A1(\bit_sel_reg[24] ),
    .A2(net259),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3445_ (.A1(_1714_),
    .A2(_1768_),
    .B(_1775_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3446_ (.A1(\bit_sel_reg[23] ),
    .A2(_1675_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3447_ (.A1(_1717_),
    .A2(net159),
    .B(_1776_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3448_ (.A1(\bit_sel_reg[22] ),
    .A2(_1675_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3449_ (.A1(_1720_),
    .A2(_1768_),
    .B(_1777_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3450_ (.A1(\bit_sel_reg[21] ),
    .A2(_1675_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3451_ (.A1(_1723_),
    .A2(_1768_),
    .B(_1778_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3452_ (.A1(\bit_sel_reg[20] ),
    .A2(_1675_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3453_ (.A1(_1726_),
    .A2(net159),
    .B(_1779_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3454_ (.A1(\bit_sel_reg[19] ),
    .A2(net258),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3455_ (.A1(_1729_),
    .A2(net159),
    .B(_1780_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3456_ (.A1(\bit_sel_reg[18] ),
    .A2(net258),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3457_ (.A1(_1732_),
    .A2(net159),
    .B(_1781_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3458_ (.A1(\bit_sel_reg[17] ),
    .A2(_1675_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3459_ (.A1(_1735_),
    .A2(net159),
    .B(_1782_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3460_ (.A1(\bit_sel_reg[16] ),
    .A2(net258),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3461_ (.A1(_1738_),
    .A2(net159),
    .B(_1783_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3462_ (.A1(\bit_sel_reg[15] ),
    .A2(_1675_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3463_ (.A1(_1740_),
    .A2(net159),
    .B(_1784_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3464_ (.A1(net5),
    .A2(_1691_),
    .A3(_1768_),
    .B1(_1676_),
    .B2(_1328_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3465_ (.A1(net5),
    .A2(_1697_),
    .A3(_1768_),
    .B1(_1676_),
    .B2(_1329_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3466_ (.A1(\bit_sel_reg[12] ),
    .A2(net259),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3467_ (.A1(_1742_),
    .A2(_1768_),
    .B(_1785_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3468_ (.A1(\bit_sel_reg[11] ),
    .A2(net258),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3469_ (.A1(_1744_),
    .A2(net159),
    .B(_1786_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3470_ (.A1(\bit_sel_reg[10] ),
    .A2(net259),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3471_ (.A1(_1746_),
    .A2(net159),
    .B(_1787_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3472_ (.A1(\bit_sel_reg[9] ),
    .A2(net258),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3473_ (.A1(_1748_),
    .A2(net159),
    .B(_1788_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3474_ (.A1(\bit_sel_reg[8] ),
    .A2(net259),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3475_ (.A1(_1750_),
    .A2(_1768_),
    .B(_1789_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3476_ (.A1(\bit_sel_reg[7] ),
    .A2(_1675_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3477_ (.A1(_1752_),
    .A2(net159),
    .B(_1790_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3478_ (.A1(\bit_sel_reg[6] ),
    .A2(_1675_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3479_ (.A1(_1754_),
    .A2(_1768_),
    .B(_1791_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3480_ (.A1(\bit_sel_reg[5] ),
    .A2(_1675_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3481_ (.A1(_1756_),
    .A2(_1768_),
    .B(_1792_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3482_ (.A1(\bit_sel_reg[4] ),
    .A2(_1675_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3483_ (.A1(_1758_),
    .A2(net159),
    .B(_1793_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3484_ (.A1(\bit_sel_reg[3] ),
    .A2(net258),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3485_ (.A1(_1760_),
    .A2(net159),
    .B(_1794_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3486_ (.A1(\bit_sel_reg[2] ),
    .A2(net258),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3487_ (.A1(_1762_),
    .A2(net159),
    .B(_1795_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3488_ (.A1(\bit_sel_reg[1] ),
    .A2(_1675_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3489_ (.A1(_1764_),
    .A2(net159),
    .B(_1796_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3490_ (.A1(\bit_sel_reg[0] ),
    .A2(net258),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3491_ (.A1(_1766_),
    .A2(net159),
    .B(_1797_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3492_ (.A1(\state[0] ),
    .A2(_1683_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3493_ (.A1(net51),
    .A2(_1363_),
    .A3(_1364_),
    .A4(_1682_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3494_ (.A1(\state[3] ),
    .A2(_1363_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3495_ (.A1(_1799_),
    .A2(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3496_ (.A1(net167),
    .A2(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3497_ (.A1(_1384_),
    .A2(_1801_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3498_ (.A1(\counter[8] ),
    .A2(_1381_),
    .A3(_1803_),
    .B(\counter[9] ),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3499_ (.A1(\state[3] ),
    .A2(_1799_),
    .B(_1804_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3500_ (.A1(_1309_),
    .A2(_1380_),
    .B(_1802_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3501_ (.A1(_1447_),
    .A2(_1801_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3502_ (.A1(_1330_),
    .A2(_1381_),
    .A3(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3503_ (.A1(_1330_),
    .A2(_1805_),
    .B(_1807_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3504_ (.A1(\counter[6] ),
    .A2(_1378_),
    .A3(_1803_),
    .B(\counter[7] ),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3505_ (.A1(_1805_),
    .A2(_1808_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3506_ (.A1(_1331_),
    .A2(_1378_),
    .A3(_1806_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3507_ (.A1(_1309_),
    .A2(_1377_),
    .B(_1802_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3508_ (.A1(_1331_),
    .A2(_1810_),
    .B(_1809_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3509_ (.A1(_1376_),
    .A2(_1803_),
    .B(\counter[5] ),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(_1810_),
    .A2(_1811_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3511_ (.A1(\state[3] ),
    .A2(_1375_),
    .B(_1803_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3512_ (.A1(_1376_),
    .A2(_1806_),
    .B1(_1812_),
    .B2(_1333_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3513_ (.A1(_1373_),
    .A2(_1802_),
    .B(_1334_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3514_ (.A1(_1812_),
    .A2(_1813_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3515_ (.A1(\counter[2] ),
    .A2(_1372_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3516_ (.A1(\counter[2] ),
    .A2(_1803_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3517_ (.A1(_1806_),
    .A2(_1814_),
    .B(_1815_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3518_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3519_ (.A1(\counter[1] ),
    .A2(_1803_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3520_ (.A1(_1806_),
    .A2(_1816_),
    .B(_1817_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3521_ (.A1(\counter[0] ),
    .A2(_1803_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3522_ (.A1(\counter[0] ),
    .A2(_1806_),
    .B(_1818_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3523_ (.A1(\state[3] ),
    .A2(_1363_),
    .B(net51),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3524_ (.A1(\state[3] ),
    .A2(_1335_),
    .B(_1385_),
    .C(_1819_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3525_ (.A1(\efuse_out[31] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[63] ),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3526_ (.A1(\efuse_out[127] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[95] ),
    .C(net9),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3527_ (.A1(_1820_),
    .A2(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3528_ (.A1(\efuse_out[191] ),
    .A2(net267),
    .B(net348),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3529_ (.A1(\efuse_out[159] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[255] ),
    .C1(net277),
    .C2(\efuse_out[223] ),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3530_ (.A1(_1823_),
    .A2(_1824_),
    .B(net361),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3531_ (.A1(\efuse_out[383] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[351] ),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3532_ (.A1(\efuse_out[287] ),
    .A2(net343),
    .B1(net367),
    .B2(\efuse_out[319] ),
    .C(net355),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3533_ (.A1(_1826_),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3534_ (.A1(\efuse_out[511] ),
    .A2(net301),
    .B(net350),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3535_ (.A1(\efuse_out[415] ),
    .A2(net341),
    .B1(net273),
    .B2(\efuse_out[479] ),
    .C1(net264),
    .C2(\efuse_out[447] ),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3536_ (.A1(_1829_),
    .A2(_1830_),
    .B(net352),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3537_ (.A1(_1822_),
    .A2(_1825_),
    .B1(_1828_),
    .B2(_1831_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3538_ (.A1(net76),
    .A2(net283),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3539_ (.A1(net283),
    .A2(_1832_),
    .B(_1833_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3540_ (.A1(\efuse_out[126] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[94] ),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3541_ (.A1(\efuse_out[30] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[62] ),
    .C(net9),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3542_ (.A1(_1834_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3543_ (.A1(\efuse_out[190] ),
    .A2(net267),
    .B(net348),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3544_ (.A1(\efuse_out[158] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[254] ),
    .C1(net277),
    .C2(\efuse_out[222] ),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3545_ (.A1(_1837_),
    .A2(_1838_),
    .B(net361),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3546_ (.A1(\efuse_out[350] ),
    .A2(net274),
    .B1(net367),
    .B2(\efuse_out[318] ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3547_ (.A1(\efuse_out[286] ),
    .A2(net343),
    .B1(net302),
    .B2(\efuse_out[382] ),
    .C(net355),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3548_ (.A1(\efuse_out[478] ),
    .A2(net273),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3549_ (.A1(\efuse_out[414] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[510] ),
    .C1(net264),
    .C2(\efuse_out[446] ),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3550_ (.A1(net355),
    .A2(_1842_),
    .A3(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3551_ (.A1(_1840_),
    .A2(_1841_),
    .B(net352),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3552_ (.A1(_1836_),
    .A2(_1839_),
    .B1(_1844_),
    .B2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3553_ (.A1(net283),
    .A2(net75),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3554_ (.A1(net283),
    .A2(_1846_),
    .B(_1847_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3555_ (.A1(\efuse_out[29] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[93] ),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3556_ (.A1(\efuse_out[125] ),
    .A2(net371),
    .B1(net261),
    .B2(\efuse_out[61] ),
    .C(net9),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3557_ (.A1(_1848_),
    .A2(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3558_ (.A1(\efuse_out[189] ),
    .A2(net267),
    .B(net348),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3559_ (.A1(\efuse_out[157] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[253] ),
    .C1(net277),
    .C2(\efuse_out[221] ),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3560_ (.A1(_1851_),
    .A2(_1852_),
    .B(net361),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3561_ (.A1(\efuse_out[285] ),
    .A2(net343),
    .B1(net302),
    .B2(\efuse_out[381] ),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3562_ (.A1(\efuse_out[349] ),
    .A2(net274),
    .B1(net367),
    .B2(\efuse_out[317] ),
    .C(net355),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3563_ (.A1(\efuse_out[445] ),
    .A2(net264),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3564_ (.A1(\efuse_out[413] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[509] ),
    .C1(net273),
    .C2(\efuse_out[477] ),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3565_ (.A1(net355),
    .A2(_1856_),
    .A3(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3566_ (.A1(_1854_),
    .A2(_1855_),
    .B(_1365_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3567_ (.A1(_1850_),
    .A2(_1853_),
    .B1(_1858_),
    .B2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3568_ (.A1(net283),
    .A2(net73),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3569_ (.A1(net283),
    .A2(_1860_),
    .B(_1861_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3570_ (.A1(\efuse_out[28] ),
    .A2(net369),
    .B1(net261),
    .B2(\efuse_out[60] ),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3571_ (.A1(\efuse_out[124] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[92] ),
    .C(net9),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3572_ (.A1(_1862_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3573_ (.A1(\efuse_out[252] ),
    .A2(net303),
    .B(net348),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3574_ (.A1(\efuse_out[156] ),
    .A2(net344),
    .B1(net277),
    .B2(\efuse_out[220] ),
    .C1(net267),
    .C2(\efuse_out[188] ),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3575_ (.A1(_1865_),
    .A2(_1866_),
    .B(net361),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3576_ (.A1(\efuse_out[380] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[348] ),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3577_ (.A1(\efuse_out[284] ),
    .A2(net343),
    .B1(net367),
    .B2(\efuse_out[316] ),
    .C(net355),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3578_ (.A1(_1868_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3579_ (.A1(\efuse_out[444] ),
    .A2(net264),
    .B(net350),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3580_ (.A1(\efuse_out[412] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[508] ),
    .C1(net273),
    .C2(\efuse_out[476] ),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3581_ (.A1(_1871_),
    .A2(_1872_),
    .B(net352),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3582_ (.A1(net158),
    .A2(_1867_),
    .B1(_1870_),
    .B2(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3583_ (.A1(net284),
    .A2(net72),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3584_ (.A1(net284),
    .A2(_1874_),
    .B(_1875_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3585_ (.A1(\efuse_out[411] ),
    .A2(net341),
    .B1(net264),
    .B2(\efuse_out[443] ),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3586_ (.A1(\efuse_out[507] ),
    .A2(net301),
    .B1(net273),
    .B2(\efuse_out[475] ),
    .C(net350),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3587_ (.A1(_1876_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3588_ (.A1(\efuse_out[283] ),
    .A2(net343),
    .B(net355),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3589_ (.A1(\efuse_out[379] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[347] ),
    .C1(\efuse_out[315] ),
    .C2(net367),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3590_ (.A1(_1879_),
    .A2(_1880_),
    .B(net352),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3591_ (.A1(\efuse_out[91] ),
    .A2(net275),
    .B1(net261),
    .B2(\efuse_out[59] ),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3592_ (.A1(\efuse_out[27] ),
    .A2(net346),
    .B1(net371),
    .B2(\efuse_out[123] ),
    .C(net355),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3593_ (.A1(\efuse_out[187] ),
    .A2(net267),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3594_ (.A1(\efuse_out[155] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[251] ),
    .C1(net277),
    .C2(\efuse_out[219] ),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3595_ (.A1(net355),
    .A2(_1884_),
    .A3(_1885_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3596_ (.A1(_1882_),
    .A2(_1883_),
    .B(net10),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3597_ (.A1(_1878_),
    .A2(_1881_),
    .B1(_1886_),
    .B2(net156),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3598_ (.A1(net283),
    .A2(net71),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3599_ (.A1(net283),
    .A2(_1888_),
    .B(_1889_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3600_ (.A1(\efuse_out[122] ),
    .A2(net371),
    .B1(net261),
    .B2(\efuse_out[58] ),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3601_ (.A1(\efuse_out[26] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[90] ),
    .C(net9),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3602_ (.A1(\efuse_out[186] ),
    .A2(net267),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3603_ (.A1(\efuse_out[154] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[250] ),
    .C1(net277),
    .C2(\efuse_out[218] ),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3604_ (.A1(net355),
    .A2(_1892_),
    .A3(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3605_ (.A1(_1890_),
    .A2(_1891_),
    .B(net10),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3606_ (.A1(\efuse_out[282] ),
    .A2(net343),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3607_ (.A1(\efuse_out[378] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[346] ),
    .C1(\efuse_out[314] ),
    .C2(net367),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3608_ (.A1(_1367_),
    .A2(_1896_),
    .A3(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3609_ (.A1(\efuse_out[410] ),
    .A2(net341),
    .B1(net273),
    .B2(\efuse_out[474] ),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3610_ (.A1(\efuse_out[506] ),
    .A2(net301),
    .B1(net264),
    .B2(\efuse_out[442] ),
    .C(net350),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3611_ (.A1(_1899_),
    .A2(_1900_),
    .B(net352),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3612_ (.A1(_1894_),
    .A2(net154),
    .B1(_1898_),
    .B2(net153),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3613_ (.A1(net284),
    .A2(net70),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3614_ (.A1(net284),
    .A2(_1902_),
    .B(_1903_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3615_ (.A1(\efuse_out[121] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[89] ),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3616_ (.A1(\efuse_out[25] ),
    .A2(net369),
    .B1(net261),
    .B2(\efuse_out[57] ),
    .C(net9),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3617_ (.A1(_1904_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3618_ (.A1(\efuse_out[217] ),
    .A2(net277),
    .B(net348),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3619_ (.A1(\efuse_out[153] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[249] ),
    .C1(net267),
    .C2(\efuse_out[185] ),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3620_ (.A1(_1907_),
    .A2(_1908_),
    .B(net360),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3621_ (.A1(\efuse_out[281] ),
    .A2(net343),
    .B1(net274),
    .B2(\efuse_out[345] ),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3622_ (.A1(\efuse_out[377] ),
    .A2(net302),
    .B1(net367),
    .B2(\efuse_out[313] ),
    .C(net355),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3623_ (.A1(_1910_),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3624_ (.A1(\efuse_out[409] ),
    .A2(net341),
    .B(net350),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3625_ (.A1(\efuse_out[505] ),
    .A2(net301),
    .B1(net273),
    .B2(\efuse_out[473] ),
    .C1(\efuse_out[441] ),
    .C2(net264),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3626_ (.A1(_1913_),
    .A2(_1914_),
    .B(net352),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3627_ (.A1(_1906_),
    .A2(_1909_),
    .B1(_1912_),
    .B2(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3628_ (.A1(net284),
    .A2(net69),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3629_ (.A1(net284),
    .A2(_1916_),
    .B(_1917_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3630_ (.A1(\efuse_out[24] ),
    .A2(net346),
    .B1(net372),
    .B2(\efuse_out[120] ),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3631_ (.A1(\efuse_out[88] ),
    .A2(net275),
    .B1(net261),
    .B2(\efuse_out[56] ),
    .C(net9),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3632_ (.A1(_1918_),
    .A2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3633_ (.A1(\efuse_out[216] ),
    .A2(net277),
    .B(net348),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3634_ (.A1(\efuse_out[152] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[248] ),
    .C1(net267),
    .C2(\efuse_out[184] ),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3635_ (.A1(_1921_),
    .A2(_1922_),
    .B(net360),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3636_ (.A1(\efuse_out[376] ),
    .A2(net302),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3637_ (.A1(_1366_),
    .A2(net7),
    .A3(\efuse_out[312] ),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3638_ (.A1(net8),
    .A2(_1368_),
    .A3(\efuse_out[344] ),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3639_ (.A1(\efuse_out[280] ),
    .A2(net343),
    .B(net355),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3640_ (.A1(_1924_),
    .A2(_1925_),
    .A3(_1926_),
    .A4(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3641_ (.A1(\efuse_out[472] ),
    .A2(net273),
    .B1(net264),
    .B2(\efuse_out[440] ),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3642_ (.A1(\efuse_out[408] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[504] ),
    .C(net350),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3643_ (.A1(_1929_),
    .A2(_1930_),
    .B(_1928_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3644_ (.A1(_1920_),
    .A2(_1923_),
    .B1(net152),
    .B2(net361),
    .C(net281),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3645_ (.A1(net283),
    .A2(net68),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3646_ (.A1(net98),
    .A2(_1933_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3647_ (.A1(\efuse_out[87] ),
    .A2(net275),
    .B1(net261),
    .B2(\efuse_out[55] ),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3648_ (.A1(\efuse_out[23] ),
    .A2(net346),
    .B1(net371),
    .B2(\efuse_out[119] ),
    .C(net9),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3649_ (.A1(_1934_),
    .A2(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3650_ (.A1(\efuse_out[215] ),
    .A2(net277),
    .B(net348),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3651_ (.A1(\efuse_out[151] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[247] ),
    .C1(net267),
    .C2(\efuse_out[183] ),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3652_ (.A1(_1937_),
    .A2(_1938_),
    .B(net360),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3653_ (.A1(\efuse_out[375] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[343] ),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3654_ (.A1(\efuse_out[279] ),
    .A2(net343),
    .B1(net367),
    .B2(\efuse_out[311] ),
    .C(net355),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3655_ (.A1(\efuse_out[439] ),
    .A2(net264),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3656_ (.A1(\efuse_out[407] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[503] ),
    .C1(net273),
    .C2(\efuse_out[471] ),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3657_ (.A1(net355),
    .A2(_1942_),
    .A3(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3658_ (.A1(_1940_),
    .A2(_1941_),
    .B(_1365_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3659_ (.A1(net151),
    .A2(_1939_),
    .B1(_1944_),
    .B2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3660_ (.A1(net285),
    .A2(net67),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3661_ (.A1(net285),
    .A2(_1946_),
    .B(_1947_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3662_ (.A1(\efuse_out[118] ),
    .A2(net373),
    .B1(net261),
    .B2(\efuse_out[54] ),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3663_ (.A1(\efuse_out[22] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[86] ),
    .C(net9),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3664_ (.A1(_1948_),
    .A2(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3665_ (.A1(\efuse_out[182] ),
    .A2(net263),
    .B(net347),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3666_ (.A1(\efuse_out[150] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[246] ),
    .C1(net277),
    .C2(\efuse_out[214] ),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3667_ (.A1(_1951_),
    .A2(_1952_),
    .B(net360),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_1950_),
    .A2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3669_ (.A1(\efuse_out[278] ),
    .A2(net343),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3670_ (.A1(\efuse_out[374] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[342] ),
    .C1(\efuse_out[310] ),
    .C2(net266),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3671_ (.A1(net350),
    .A2(_1955_),
    .A3(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3672_ (.A1(\efuse_out[406] ),
    .A2(net341),
    .B1(net273),
    .B2(\efuse_out[470] ),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3673_ (.A1(\efuse_out[502] ),
    .A2(net301),
    .B1(net264),
    .B2(\efuse_out[438] ),
    .C(net350),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3674_ (.A1(_1958_),
    .A2(_1959_),
    .B(net352),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3675_ (.A1(_1957_),
    .A2(_1960_),
    .B(net279),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3676_ (.A1(net279),
    .A2(_1336_),
    .B1(_1954_),
    .B2(_1961_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3677_ (.A1(\efuse_out[21] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[53] ),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3678_ (.A1(\efuse_out[117] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[85] ),
    .C(net9),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3679_ (.A1(_1962_),
    .A2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3680_ (.A1(\efuse_out[245] ),
    .A2(net303),
    .B(net348),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3681_ (.A1(\efuse_out[149] ),
    .A2(net345),
    .B1(net277),
    .B2(\efuse_out[213] ),
    .C1(net263),
    .C2(\efuse_out[181] ),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3682_ (.A1(_1965_),
    .A2(_1966_),
    .B(net360),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3683_ (.A1(\efuse_out[373] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[341] ),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3684_ (.A1(\efuse_out[277] ),
    .A2(net343),
    .B1(net266),
    .B2(\efuse_out[309] ),
    .C(net355),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3685_ (.A1(_1968_),
    .A2(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3686_ (.A1(\efuse_out[405] ),
    .A2(net341),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3687_ (.A1(\efuse_out[501] ),
    .A2(net301),
    .B1(net273),
    .B2(\efuse_out[469] ),
    .C1(\efuse_out[437] ),
    .C2(net264),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3688_ (.A1(net355),
    .A2(_1971_),
    .A3(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3689_ (.A1(net361),
    .A2(_1970_),
    .A3(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3690_ (.A1(_1964_),
    .A2(_1967_),
    .B(net281),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3691_ (.A1(net279),
    .A2(_1337_),
    .B1(_1974_),
    .B2(net97),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3692_ (.A1(\efuse_out[500] ),
    .A2(net301),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3693_ (.A1(\efuse_out[404] ),
    .A2(net341),
    .B1(net273),
    .B2(\efuse_out[468] ),
    .C1(net264),
    .C2(\efuse_out[436] ),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3694_ (.A1(net355),
    .A2(_1976_),
    .A3(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3695_ (.A1(\efuse_out[372] ),
    .A2(net302),
    .B1(net266),
    .B2(\efuse_out[308] ),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3696_ (.A1(\efuse_out[276] ),
    .A2(net343),
    .B1(net274),
    .B2(\efuse_out[340] ),
    .C(net355),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3697_ (.A1(_1979_),
    .A2(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3698_ (.A1(net361),
    .A2(_1978_),
    .A3(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3699_ (.A1(\efuse_out[116] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[84] ),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3700_ (.A1(\efuse_out[20] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[52] ),
    .C(net9),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3701_ (.A1(_1983_),
    .A2(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3702_ (.A1(\efuse_out[244] ),
    .A2(net303),
    .B(net348),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3703_ (.A1(\efuse_out[148] ),
    .A2(net345),
    .B1(net277),
    .B2(\efuse_out[212] ),
    .C1(net262),
    .C2(\efuse_out[180] ),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3704_ (.A1(_1986_),
    .A2(_1987_),
    .B(net360),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3705_ (.A1(_1985_),
    .A2(_1988_),
    .B(net281),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3706_ (.A1(net279),
    .A2(_1338_),
    .B1(_1982_),
    .B2(net96),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3707_ (.A1(\efuse_out[19] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[83] ),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3708_ (.A1(\efuse_out[115] ),
    .A2(net373),
    .B1(net263),
    .B2(\efuse_out[51] ),
    .C(net9),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3709_ (.A1(_1990_),
    .A2(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3710_ (.A1(\efuse_out[179] ),
    .A2(net262),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3711_ (.A1(\efuse_out[147] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[243] ),
    .C1(net276),
    .C2(\efuse_out[211] ),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3712_ (.A1(net9),
    .A2(_1993_),
    .A3(_1994_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3713_ (.A1(net354),
    .A2(_1992_),
    .A3(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3714_ (.A1(\efuse_out[339] ),
    .A2(net274),
    .B(net355),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3715_ (.A1(\efuse_out[275] ),
    .A2(net343),
    .B1(net302),
    .B2(\efuse_out[371] ),
    .C1(net266),
    .C2(\efuse_out[307] ),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3716_ (.A1(\efuse_out[499] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[467] ),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3717_ (.A1(\efuse_out[403] ),
    .A2(net341),
    .B1(net264),
    .B2(\efuse_out[435] ),
    .C(net350),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3718_ (.A1(_1999_),
    .A2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3719_ (.A1(_1997_),
    .A2(_1998_),
    .B(net352),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3720_ (.A1(_2001_),
    .A2(_2002_),
    .B(net279),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3721_ (.A1(net279),
    .A2(_1339_),
    .B1(_1996_),
    .B2(_2003_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3722_ (.A1(\efuse_out[114] ),
    .A2(net374),
    .B1(net263),
    .B2(\efuse_out[50] ),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3723_ (.A1(\efuse_out[18] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[82] ),
    .C(net9),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3724_ (.A1(_2004_),
    .A2(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3725_ (.A1(\efuse_out[242] ),
    .A2(net303),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3726_ (.A1(\efuse_out[146] ),
    .A2(net345),
    .B1(net277),
    .B2(\efuse_out[210] ),
    .C1(net262),
    .C2(\efuse_out[178] ),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3727_ (.A1(net9),
    .A2(_2007_),
    .A3(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3728_ (.A1(net354),
    .A2(_2006_),
    .A3(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(\efuse_out[370] ),
    .A2(net302),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3730_ (.A1(\efuse_out[274] ),
    .A2(net343),
    .B1(net364),
    .B2(\efuse_out[338] ),
    .C1(net265),
    .C2(\efuse_out[306] ),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3731_ (.A1(net350),
    .A2(_2011_),
    .A3(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3732_ (.A1(\efuse_out[402] ),
    .A2(net341),
    .B1(net272),
    .B2(\efuse_out[466] ),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3733_ (.A1(\efuse_out[498] ),
    .A2(net301),
    .B1(net264),
    .B2(\efuse_out[434] ),
    .C(net349),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3734_ (.A1(_2014_),
    .A2(_2015_),
    .B(net352),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3735_ (.A1(_2013_),
    .A2(_2016_),
    .B(net279),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3736_ (.A1(net279),
    .A2(_1340_),
    .B1(_2010_),
    .B2(_2017_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3737_ (.A1(\efuse_out[113] ),
    .A2(net374),
    .B1(net263),
    .B2(\efuse_out[49] ),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3738_ (.A1(\efuse_out[17] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[81] ),
    .C(net9),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3739_ (.A1(_2018_),
    .A2(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3740_ (.A1(\efuse_out[177] ),
    .A2(net262),
    .B(net347),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3741_ (.A1(\efuse_out[145] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[241] ),
    .C1(net276),
    .C2(\efuse_out[209] ),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3742_ (.A1(_2021_),
    .A2(_2022_),
    .B(net360),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3743_ (.A1(\efuse_out[369] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[337] ),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3744_ (.A1(\efuse_out[273] ),
    .A2(net343),
    .B1(net266),
    .B2(\efuse_out[305] ),
    .C(net355),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3745_ (.A1(\efuse_out[465] ),
    .A2(net272),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3746_ (.A1(\efuse_out[401] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[497] ),
    .C1(net264),
    .C2(\efuse_out[433] ),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3747_ (.A1(net355),
    .A2(_2026_),
    .A3(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3748_ (.A1(_2024_),
    .A2(_2025_),
    .B(net351),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3749_ (.A1(_2020_),
    .A2(_2023_),
    .B1(_2028_),
    .B2(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3750_ (.A1(net283),
    .A2(net60),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3751_ (.A1(net284),
    .A2(_2030_),
    .B(_2031_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3752_ (.A1(\efuse_out[400] ),
    .A2(net341),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3753_ (.A1(\efuse_out[496] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[464] ),
    .C1(\efuse_out[432] ),
    .C2(net264),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3754_ (.A1(net355),
    .A2(_2032_),
    .A3(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3755_ (.A1(\efuse_out[272] ),
    .A2(net343),
    .B1(net364),
    .B2(\efuse_out[336] ),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3756_ (.A1(\efuse_out[368] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[304] ),
    .C(net355),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3757_ (.A1(_2035_),
    .A2(_2036_),
    .B(net351),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3758_ (.A1(\efuse_out[16] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[80] ),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3759_ (.A1(\efuse_out[112] ),
    .A2(net374),
    .B1(net263),
    .B2(\efuse_out[48] ),
    .C(net9),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3760_ (.A1(_2038_),
    .A2(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3761_ (.A1(\efuse_out[144] ),
    .A2(net345),
    .B(net347),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3762_ (.A1(\efuse_out[240] ),
    .A2(net303),
    .B1(net276),
    .B2(\efuse_out[208] ),
    .C1(\efuse_out[176] ),
    .C2(net267),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3763_ (.A1(_2041_),
    .A2(_2042_),
    .B(net360),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3764_ (.A1(_2034_),
    .A2(_2037_),
    .B1(_2040_),
    .B2(_2043_),
    .C(net280),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3765_ (.A1(net284),
    .A2(net59),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3766_ (.A1(net95),
    .A2(_2045_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3767_ (.A1(\efuse_out[79] ),
    .A2(net275),
    .B1(net263),
    .B2(\efuse_out[47] ),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3768_ (.A1(\efuse_out[15] ),
    .A2(net346),
    .B1(net374),
    .B2(\efuse_out[111] ),
    .C(net9),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3769_ (.A1(_2046_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3770_ (.A1(\efuse_out[207] ),
    .A2(net277),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3771_ (.A1(\efuse_out[143] ),
    .A2(net345),
    .B1(net303),
    .B2(\efuse_out[239] ),
    .C1(net262),
    .C2(\efuse_out[175] ),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3772_ (.A1(net9),
    .A2(_2049_),
    .A3(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3773_ (.A1(net354),
    .A2(_2048_),
    .A3(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3774_ (.A1(\efuse_out[271] ),
    .A2(net342),
    .B1(net274),
    .B2(\efuse_out[335] ),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3775_ (.A1(\efuse_out[367] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[303] ),
    .C(net355),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3776_ (.A1(_2053_),
    .A2(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3777_ (.A1(\efuse_out[495] ),
    .A2(net301),
    .B(net349),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3778_ (.A1(\efuse_out[399] ),
    .A2(net341),
    .B1(net272),
    .B2(\efuse_out[463] ),
    .C1(net264),
    .C2(\efuse_out[431] ),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3779_ (.A1(_2056_),
    .A2(_2057_),
    .B(net352),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3780_ (.A1(_2055_),
    .A2(_2058_),
    .B(net279),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3781_ (.A1(net279),
    .A2(_1341_),
    .B1(_2052_),
    .B2(_2059_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3782_ (.A1(\efuse_out[14] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[46] ),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3783_ (.A1(\efuse_out[110] ),
    .A2(net374),
    .B1(net275),
    .B2(\efuse_out[78] ),
    .C(net9),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3784_ (.A1(_2060_),
    .A2(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3785_ (.A1(\efuse_out[174] ),
    .A2(net262),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3786_ (.A1(\efuse_out[142] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[238] ),
    .C1(net276),
    .C2(\efuse_out[206] ),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3787_ (.A1(net9),
    .A2(_2063_),
    .A3(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3788_ (.A1(net353),
    .A2(_2062_),
    .A3(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3789_ (.A1(\efuse_out[334] ),
    .A2(net274),
    .B(net355),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3790_ (.A1(\efuse_out[270] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[366] ),
    .C1(net265),
    .C2(\efuse_out[302] ),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3791_ (.A1(\efuse_out[494] ),
    .A2(net301),
    .B1(net264),
    .B2(\efuse_out[430] ),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3792_ (.A1(\efuse_out[398] ),
    .A2(net341),
    .B1(net272),
    .B2(\efuse_out[462] ),
    .C(net349),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3793_ (.A1(_2069_),
    .A2(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3794_ (.A1(_2067_),
    .A2(_2068_),
    .B(net351),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3795_ (.A1(_2071_),
    .A2(_2072_),
    .B(net279),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3796_ (.A1(net279),
    .A2(_1342_),
    .B1(_2066_),
    .B2(_2073_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3797_ (.A1(\efuse_out[461] ),
    .A2(net272),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3798_ (.A1(\efuse_out[397] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[493] ),
    .C1(net264),
    .C2(\efuse_out[429] ),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3799_ (.A1(net355),
    .A2(_2074_),
    .A3(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3800_ (.A1(\efuse_out[269] ),
    .A2(net342),
    .B1(net274),
    .B2(\efuse_out[333] ),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3801_ (.A1(\efuse_out[365] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[301] ),
    .C(net355),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(_2077_),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3803_ (.A1(net361),
    .A2(_2076_),
    .A3(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3804_ (.A1(\efuse_out[13] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[45] ),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3805_ (.A1(\efuse_out[109] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[77] ),
    .C(net9),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3806_ (.A1(_2081_),
    .A2(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3807_ (.A1(\efuse_out[205] ),
    .A2(net277),
    .B(net347),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3808_ (.A1(\efuse_out[141] ),
    .A2(net345),
    .B1(net303),
    .B2(\efuse_out[237] ),
    .C1(net262),
    .C2(\efuse_out[173] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3809_ (.A1(_2084_),
    .A2(_2085_),
    .B(net360),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3810_ (.A1(_2083_),
    .A2(_2086_),
    .B(_1335_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3811_ (.A1(net279),
    .A2(_1343_),
    .B1(_2080_),
    .B2(net94),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3812_ (.A1(\efuse_out[396] ),
    .A2(net341),
    .B1(net264),
    .B2(\efuse_out[428] ),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3813_ (.A1(\efuse_out[492] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[460] ),
    .C(net349),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3814_ (.A1(_2088_),
    .A2(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3815_ (.A1(\efuse_out[300] ),
    .A2(net265),
    .B(net355),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3816_ (.A1(\efuse_out[268] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[364] ),
    .C1(net274),
    .C2(\efuse_out[332] ),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3817_ (.A1(_2091_),
    .A2(_2092_),
    .B(net351),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3818_ (.A1(\efuse_out[12] ),
    .A2(net346),
    .B1(net371),
    .B2(\efuse_out[108] ),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3819_ (.A1(\efuse_out[76] ),
    .A2(net275),
    .B1(net263),
    .B2(\efuse_out[44] ),
    .C(net9),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3820_ (.A1(\efuse_out[140] ),
    .A2(net344),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3821_ (.A1(\efuse_out[236] ),
    .A2(net303),
    .B1(net276),
    .B2(\efuse_out[204] ),
    .C1(\efuse_out[172] ),
    .C2(net267),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3822_ (.A1(net9),
    .A2(_2096_),
    .A3(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3823_ (.A1(_2094_),
    .A2(_2095_),
    .B(net10),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3824_ (.A1(_2090_),
    .A2(_2093_),
    .B1(_2098_),
    .B2(net149),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3825_ (.A1(net283),
    .A2(net55),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3826_ (.A1(net283),
    .A2(net93),
    .B(_2101_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3827_ (.A1(\efuse_out[11] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[43] ),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3828_ (.A1(\efuse_out[107] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[75] ),
    .C(net9),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3829_ (.A1(_2102_),
    .A2(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3830_ (.A1(\efuse_out[203] ),
    .A2(net277),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3831_ (.A1(\efuse_out[139] ),
    .A2(net345),
    .B1(net303),
    .B2(\efuse_out[235] ),
    .C1(net262),
    .C2(\efuse_out[171] ),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3832_ (.A1(net9),
    .A2(_2105_),
    .A3(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3833_ (.A1(net353),
    .A2(_2104_),
    .A3(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3834_ (.A1(\efuse_out[267] ),
    .A2(net342),
    .B1(net274),
    .B2(\efuse_out[331] ),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3835_ (.A1(\efuse_out[363] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[299] ),
    .C(net355),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(\efuse_out[459] ),
    .A2(net272),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3837_ (.A1(\efuse_out[395] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[491] ),
    .C1(net264),
    .C2(\efuse_out[427] ),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3838_ (.A1(net355),
    .A2(_2111_),
    .A3(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3839_ (.A1(_2109_),
    .A2(_2110_),
    .B(net351),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3840_ (.A1(_2113_),
    .A2(_2114_),
    .B(net278),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3841_ (.A1(net278),
    .A2(_1344_),
    .B1(_2108_),
    .B2(_2115_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(\efuse_out[394] ),
    .A2(net341),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3843_ (.A1(\efuse_out[490] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[458] ),
    .C1(\efuse_out[426] ),
    .C2(net264),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3844_ (.A1(net355),
    .A2(_2116_),
    .A3(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3845_ (.A1(\efuse_out[266] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[362] ),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3846_ (.A1(\efuse_out[330] ),
    .A2(net364),
    .B1(net265),
    .B2(\efuse_out[298] ),
    .C(net355),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3847_ (.A1(_2119_),
    .A2(_2120_),
    .B(net351),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3848_ (.A1(\efuse_out[106] ),
    .A2(net374),
    .B1(net263),
    .B2(\efuse_out[42] ),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3849_ (.A1(\efuse_out[10] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[74] ),
    .C(net9),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3850_ (.A1(_2122_),
    .A2(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3851_ (.A1(\efuse_out[234] ),
    .A2(net303),
    .B(net348),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3852_ (.A1(\efuse_out[138] ),
    .A2(net345),
    .B1(net277),
    .B2(\efuse_out[202] ),
    .C1(net262),
    .C2(\efuse_out[170] ),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3853_ (.A1(_2125_),
    .A2(_2126_),
    .B(net360),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3854_ (.A1(_2118_),
    .A2(_2121_),
    .B1(_2124_),
    .B2(_2127_),
    .C(net278),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3855_ (.A1(net283),
    .A2(net53),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3856_ (.A1(net91),
    .A2(_2129_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3857_ (.A1(\efuse_out[9] ),
    .A2(net346),
    .B1(net371),
    .B2(\efuse_out[105] ),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3858_ (.A1(\efuse_out[73] ),
    .A2(net275),
    .B1(net263),
    .B2(\efuse_out[41] ),
    .C(net9),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3859_ (.A1(_2130_),
    .A2(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3860_ (.A1(\efuse_out[169] ),
    .A2(net262),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3861_ (.A1(\efuse_out[137] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[233] ),
    .C1(net276),
    .C2(\efuse_out[201] ),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3862_ (.A1(net9),
    .A2(_2133_),
    .A3(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3863_ (.A1(net353),
    .A2(_2132_),
    .A3(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3864_ (.A1(\efuse_out[265] ),
    .A2(net342),
    .B1(net274),
    .B2(\efuse_out[329] ),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3865_ (.A1(\efuse_out[361] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[297] ),
    .C(net355),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3866_ (.A1(\efuse_out[393] ),
    .A2(net341),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3867_ (.A1(\efuse_out[489] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[457] ),
    .C1(\efuse_out[425] ),
    .C2(net264),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3868_ (.A1(net355),
    .A2(_2139_),
    .A3(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3869_ (.A1(_2137_),
    .A2(_2138_),
    .B(net351),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3870_ (.A1(_2141_),
    .A2(_2142_),
    .B(net278),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3871_ (.A1(net278),
    .A2(_1345_),
    .B1(_2136_),
    .B2(_2143_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3872_ (.A1(\efuse_out[456] ),
    .A2(net272),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3873_ (.A1(\efuse_out[392] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[488] ),
    .C1(net264),
    .C2(\efuse_out[424] ),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3874_ (.A1(net355),
    .A2(_2144_),
    .A3(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3875_ (.A1(\efuse_out[360] ),
    .A2(net302),
    .B1(net265),
    .B2(\efuse_out[296] ),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3876_ (.A1(\efuse_out[264] ),
    .A2(net342),
    .B1(net274),
    .B2(\efuse_out[328] ),
    .C(net355),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3877_ (.A1(_2147_),
    .A2(_2148_),
    .B(net351),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3878_ (.A1(\efuse_out[8] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[40] ),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3879_ (.A1(\efuse_out[104] ),
    .A2(net375),
    .B1(net275),
    .B2(\efuse_out[72] ),
    .C(net9),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3880_ (.A1(_2150_),
    .A2(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3881_ (.A1(\efuse_out[168] ),
    .A2(net262),
    .B(net347),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3882_ (.A1(\efuse_out[136] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[232] ),
    .C1(net276),
    .C2(\efuse_out[200] ),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3883_ (.A1(_2153_),
    .A2(_2154_),
    .B(net360),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3884_ (.A1(_2146_),
    .A2(_2149_),
    .B1(_2152_),
    .B2(_2155_),
    .C(net278),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3885_ (.A1(net283),
    .A2(net82),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3886_ (.A1(net90),
    .A2(_2157_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3887_ (.A1(\efuse_out[7] ),
    .A2(net370),
    .B1(net261),
    .B2(\efuse_out[39] ),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3888_ (.A1(\efuse_out[103] ),
    .A2(net375),
    .B1(net275),
    .B2(\efuse_out[71] ),
    .C(net9),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3889_ (.A1(_2158_),
    .A2(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3890_ (.A1(\efuse_out[199] ),
    .A2(net276),
    .B(net348),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3891_ (.A1(\efuse_out[135] ),
    .A2(net345),
    .B1(net303),
    .B2(\efuse_out[231] ),
    .C1(net262),
    .C2(\efuse_out[167] ),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3892_ (.A1(_2161_),
    .A2(_2162_),
    .B(net360),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3893_ (.A1(\efuse_out[359] ),
    .A2(net302),
    .B1(net274),
    .B2(\efuse_out[327] ),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3894_ (.A1(\efuse_out[263] ),
    .A2(net342),
    .B1(net265),
    .B2(\efuse_out[295] ),
    .C(net9),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3895_ (.A1(\efuse_out[391] ),
    .A2(net341),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3896_ (.A1(\efuse_out[487] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[455] ),
    .C1(\efuse_out[423] ),
    .C2(net264),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3897_ (.A1(net355),
    .A2(_2166_),
    .A3(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3898_ (.A1(_2164_),
    .A2(_2165_),
    .B(net351),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3899_ (.A1(_2160_),
    .A2(_2163_),
    .B1(_2168_),
    .B2(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3900_ (.A1(net283),
    .A2(net81),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3901_ (.A1(net283),
    .A2(net89),
    .B(_2171_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3902_ (.A1(\efuse_out[102] ),
    .A2(net371),
    .B1(net263),
    .B2(\efuse_out[38] ),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3903_ (.A1(\efuse_out[6] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[70] ),
    .C(net9),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3904_ (.A1(_2172_),
    .A2(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3905_ (.A1(\efuse_out[166] ),
    .A2(net262),
    .B(net347),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3906_ (.A1(\efuse_out[134] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[230] ),
    .C1(net276),
    .C2(\efuse_out[198] ),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3907_ (.A1(_2175_),
    .A2(_2176_),
    .B(net360),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3908_ (.A1(\efuse_out[326] ),
    .A2(net365),
    .B1(net265),
    .B2(\efuse_out[294] ),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3909_ (.A1(\efuse_out[262] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[358] ),
    .C(net355),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3910_ (.A1(\efuse_out[390] ),
    .A2(net341),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3911_ (.A1(\efuse_out[486] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[454] ),
    .C1(\efuse_out[422] ),
    .C2(net264),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3912_ (.A1(net355),
    .A2(_2180_),
    .A3(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3913_ (.A1(_2178_),
    .A2(_2179_),
    .B(net351),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3914_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2182_),
    .B2(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3915_ (.A1(net283),
    .A2(net80),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3916_ (.A1(net283),
    .A2(net88),
    .B(_2185_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3917_ (.A1(\efuse_out[485] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[453] ),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3918_ (.A1(\efuse_out[389] ),
    .A2(net341),
    .B1(net264),
    .B2(\efuse_out[421] ),
    .C(net349),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3919_ (.A1(_2186_),
    .A2(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3920_ (.A1(\efuse_out[325] ),
    .A2(net365),
    .B(net355),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3921_ (.A1(\efuse_out[261] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[357] ),
    .C1(net265),
    .C2(\efuse_out[293] ),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3922_ (.A1(_2189_),
    .A2(_2190_),
    .B(net351),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3923_ (.A1(\efuse_out[5] ),
    .A2(net368),
    .B1(net261),
    .B2(\efuse_out[37] ),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3924_ (.A1(\efuse_out[101] ),
    .A2(net371),
    .B1(net275),
    .B2(\efuse_out[69] ),
    .C(net9),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3925_ (.A1(\efuse_out[165] ),
    .A2(net262),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3926_ (.A1(\efuse_out[133] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[229] ),
    .C1(net276),
    .C2(\efuse_out[197] ),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3927_ (.A1(net9),
    .A2(_2194_),
    .A3(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3928_ (.A1(_2192_),
    .A2(_2193_),
    .B(net10),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3929_ (.A1(_2188_),
    .A2(_2191_),
    .B1(_2196_),
    .B2(net147),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3930_ (.A1(net284),
    .A2(net79),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3931_ (.A1(net284),
    .A2(net87),
    .B(_2199_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3932_ (.A1(\efuse_out[4] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[68] ),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3933_ (.A1(\efuse_out[100] ),
    .A2(net375),
    .B1(net263),
    .B2(\efuse_out[36] ),
    .C(net9),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(_2200_),
    .A2(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3935_ (.A1(\efuse_out[132] ),
    .A2(net345),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3936_ (.A1(\efuse_out[228] ),
    .A2(net303),
    .B1(net276),
    .B2(\efuse_out[196] ),
    .C1(\efuse_out[164] ),
    .C2(net262),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3937_ (.A1(net9),
    .A2(_2203_),
    .A3(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3938_ (.A1(net353),
    .A2(_2202_),
    .A3(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3939_ (.A1(\efuse_out[292] ),
    .A2(net265),
    .B(net355),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3940_ (.A1(\efuse_out[260] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[356] ),
    .C1(net364),
    .C2(\efuse_out[324] ),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3941_ (.A1(\efuse_out[484] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[452] ),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3942_ (.A1(\efuse_out[388] ),
    .A2(net341),
    .B1(net264),
    .B2(\efuse_out[420] ),
    .C(net349),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(_2209_),
    .A2(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3944_ (.A1(_2207_),
    .A2(_2208_),
    .B(net351),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3945_ (.A1(_2211_),
    .A2(_2212_),
    .B(net278),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3946_ (.A1(net278),
    .A2(_1346_),
    .B1(_2206_),
    .B2(_2213_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3947_ (.A1(\efuse_out[3] ),
    .A2(net370),
    .B(net9),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3948_ (.A1(\efuse_out[99] ),
    .A2(net372),
    .B1(net275),
    .B2(\efuse_out[67] ),
    .C1(\efuse_out[35] ),
    .C2(net263),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3949_ (.A1(\efuse_out[163] ),
    .A2(net262),
    .B(net347),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3950_ (.A1(\efuse_out[131] ),
    .A2(net345),
    .B1(net303),
    .B2(\efuse_out[227] ),
    .C1(net276),
    .C2(\efuse_out[195] ),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3951_ (.A1(_2214_),
    .A2(net181),
    .B1(_2216_),
    .B2(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3952_ (.A1(\efuse_out[355] ),
    .A2(net302),
    .B(net355),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3953_ (.A1(\efuse_out[259] ),
    .A2(net342),
    .B1(net365),
    .B2(\efuse_out[323] ),
    .C1(net265),
    .C2(\efuse_out[291] ),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3954_ (.A1(\efuse_out[483] ),
    .A2(net301),
    .B1(net264),
    .B2(\efuse_out[419] ),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3955_ (.A1(\efuse_out[387] ),
    .A2(net341),
    .B1(net272),
    .B2(\efuse_out[451] ),
    .C(net349),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3956_ (.A1(_2221_),
    .A2(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3957_ (.A1(_2219_),
    .A2(_2220_),
    .B(net351),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3958_ (.A1(net351),
    .A2(net146),
    .B1(_2223_),
    .B2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3959_ (.A1(net284),
    .A2(net77),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3960_ (.A1(net284),
    .A2(net86),
    .B(_2226_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3961_ (.A1(\efuse_out[66] ),
    .A2(net275),
    .B1(net263),
    .B2(\efuse_out[34] ),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3962_ (.A1(\efuse_out[2] ),
    .A2(net346),
    .B1(net375),
    .B2(\efuse_out[98] ),
    .C(net9),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3963_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3964_ (.A1(\efuse_out[162] ),
    .A2(net262),
    .B(net348),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3965_ (.A1(\efuse_out[130] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[226] ),
    .C1(net276),
    .C2(\efuse_out[194] ),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3966_ (.A1(_2230_),
    .A2(_2231_),
    .B(net360),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3967_ (.A1(\efuse_out[258] ),
    .A2(net342),
    .B1(net265),
    .B2(\efuse_out[290] ),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3968_ (.A1(\efuse_out[354] ),
    .A2(net302),
    .B1(net364),
    .B2(\efuse_out[322] ),
    .C(net355),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3969_ (.A1(\efuse_out[418] ),
    .A2(net264),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3970_ (.A1(\efuse_out[386] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[482] ),
    .C1(net272),
    .C2(\efuse_out[450] ),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3971_ (.A1(net355),
    .A2(_2235_),
    .A3(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3972_ (.A1(_2233_),
    .A2(_2234_),
    .B(net351),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3973_ (.A1(_2229_),
    .A2(_2232_),
    .B1(_2237_),
    .B2(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3974_ (.A1(net284),
    .A2(net74),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3975_ (.A1(net284),
    .A2(net85),
    .B(_2240_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3976_ (.A1(\efuse_out[1] ),
    .A2(net346),
    .B1(net275),
    .B2(\efuse_out[65] ),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3977_ (.A1(\efuse_out[97] ),
    .A2(net375),
    .B1(net263),
    .B2(\efuse_out[33] ),
    .C(net9),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3978_ (.A1(_2241_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3979_ (.A1(\efuse_out[129] ),
    .A2(net344),
    .B(net348),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3980_ (.A1(\efuse_out[225] ),
    .A2(net303),
    .B1(net276),
    .B2(\efuse_out[193] ),
    .C1(\efuse_out[161] ),
    .C2(net262),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3981_ (.A1(_2244_),
    .A2(_2245_),
    .B(net360),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3982_ (.A1(\efuse_out[321] ),
    .A2(net365),
    .B1(net265),
    .B2(\efuse_out[289] ),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3983_ (.A1(\efuse_out[257] ),
    .A2(net342),
    .B1(net302),
    .B2(\efuse_out[353] ),
    .C(net9),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3984_ (.A1(_2247_),
    .A2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3985_ (.A1(\efuse_out[385] ),
    .A2(net341),
    .B(net349),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3986_ (.A1(\efuse_out[481] ),
    .A2(net301),
    .B1(net272),
    .B2(\efuse_out[449] ),
    .C1(\efuse_out[417] ),
    .C2(net264),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3987_ (.A1(_2250_),
    .A2(_2251_),
    .B(net351),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3988_ (.A1(net145),
    .A2(_2246_),
    .B1(_2249_),
    .B2(net144),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3989_ (.A1(net284),
    .A2(net63),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3990_ (.A1(net284),
    .A2(net84),
    .B(_2254_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3991_ (.A1(\efuse_out[0] ),
    .A2(net346),
    .B1(net375),
    .B2(\efuse_out[96] ),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3992_ (.A1(\efuse_out[64] ),
    .A2(net275),
    .B1(net263),
    .B2(\efuse_out[32] ),
    .C(net9),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3993_ (.A1(_2255_),
    .A2(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(\efuse_out[160] ),
    .A2(net262),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3995_ (.A1(\efuse_out[128] ),
    .A2(net344),
    .B1(net303),
    .B2(\efuse_out[224] ),
    .C1(net276),
    .C2(\efuse_out[192] ),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3996_ (.A1(net9),
    .A2(_2258_),
    .A3(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3997_ (.A1(net353),
    .A2(_2257_),
    .A3(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3998_ (.A1(\efuse_out[256] ),
    .A2(net342),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3999_ (.A1(\efuse_out[352] ),
    .A2(net302),
    .B1(net365),
    .B2(\efuse_out[320] ),
    .C1(\efuse_out[288] ),
    .C2(net265),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4000_ (.A1(_1367_),
    .A2(_2262_),
    .A3(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4001_ (.A1(\efuse_out[384] ),
    .A2(net341),
    .B1(net301),
    .B2(\efuse_out[480] ),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4002_ (.A1(\efuse_out[448] ),
    .A2(net272),
    .B1(net264),
    .B2(\efuse_out[416] ),
    .C(net349),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4003_ (.A1(_2265_),
    .A2(_2266_),
    .B(net351),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4004_ (.A1(_2264_),
    .A2(_2267_),
    .B(net280),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4005_ (.A1(net280),
    .A2(_1347_),
    .B1(_2261_),
    .B2(_2268_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4006_ (.A1(net51),
    .A2(net50),
    .A3(_1682_),
    .B(\state[0] ),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4007_ (.A1(\state[1] ),
    .A2(_2269_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4008_ (.A1(net9),
    .A2(net303),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4009_ (.A1(net361),
    .A2(net355),
    .A3(net302),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4010_ (.I(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4011_ (.A1(net50),
    .A2(_1798_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4012_ (.A1(_1335_),
    .A2(\state[0] ),
    .B1(net50),
    .B2(_1798_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4013_ (.A1(_2273_),
    .A2(net142),
    .B(\sense_reg[15] ),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4014_ (.A1(net180),
    .A2(_2275_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4015_ (.A1(net8),
    .A2(net9),
    .A3(_1368_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4016_ (.A1(net353),
    .A2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4017_ (.A1(net361),
    .A2(net355),
    .A3(net274),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4018_ (.A1(net142),
    .A2(net179),
    .B(\sense_reg[14] ),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4019_ (.A1(net180),
    .A2(_2279_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4020_ (.A1(_1366_),
    .A2(net9),
    .A3(net7),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4021_ (.A1(net353),
    .A2(_2280_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4022_ (.A1(net361),
    .A2(net355),
    .A3(net265),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4023_ (.A1(net142),
    .A2(net178),
    .B(\sense_reg[13] ),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4024_ (.A1(net180),
    .A2(_2283_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4025_ (.A1(net352),
    .A2(net350),
    .A3(_1387_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4026_ (.A1(net361),
    .A2(net355),
    .A3(net342),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4027_ (.A1(net142),
    .A2(_2284_),
    .B(\sense_reg[12] ),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4028_ (.A1(net180),
    .A2(_2286_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4029_ (.A1(net351),
    .A2(net355),
    .A3(_1473_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4030_ (.A1(net361),
    .A2(net350),
    .A3(net302),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4031_ (.A1(net142),
    .A2(net256),
    .B(\sense_reg[11] ),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4032_ (.A1(net180),
    .A2(_2289_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4033_ (.A1(net353),
    .A2(_1531_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4034_ (.A1(net360),
    .A2(_1367_),
    .A3(net276),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4035_ (.A1(net142),
    .A2(_2290_),
    .B(\sense_reg[10] ),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4036_ (.A1(net180),
    .A2(_2292_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4037_ (.A1(net353),
    .A2(_1590_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4038_ (.A1(net360),
    .A2(_1367_),
    .A3(net267),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4039_ (.A1(net142),
    .A2(_2293_),
    .B(\sense_reg[9] ),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4040_ (.A1(net180),
    .A2(_2295_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4041_ (.A1(net360),
    .A2(net288),
    .A3(net142),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4042_ (.A1(_1348_),
    .A2(_2296_),
    .B(net180),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4043_ (.A1(net360),
    .A2(_2271_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4044_ (.A1(net353),
    .A2(net9),
    .A3(net303),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4045_ (.A1(net142),
    .A2(_2297_),
    .B(\sense_reg[7] ),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4046_ (.A1(net180),
    .A2(_2299_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4047_ (.A1(net360),
    .A2(_2276_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4048_ (.A1(net353),
    .A2(net9),
    .A3(net276),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4049_ (.A1(net143),
    .A2(_2300_),
    .B(\sense_reg[6] ),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4050_ (.A1(_2270_),
    .A2(_2302_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4051_ (.A1(net360),
    .A2(_2280_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4052_ (.A1(net353),
    .A2(net9),
    .A3(net262),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4053_ (.A1(net143),
    .A2(_2303_),
    .B(\sense_reg[5] ),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4054_ (.A1(_2270_),
    .A2(_2305_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4055_ (.A1(_1388_),
    .A2(net143),
    .B(\sense_reg[4] ),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4056_ (.A1(_2270_),
    .A2(_2306_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4057_ (.A1(_1474_),
    .A2(net143),
    .B(\sense_reg[3] ),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4058_ (.A1(_2270_),
    .A2(_2307_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4059_ (.A1(_1532_),
    .A2(net143),
    .B(\sense_reg[2] ),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4060_ (.A1(_2270_),
    .A2(_2308_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4061_ (.A1(_1591_),
    .A2(net143),
    .B(\sense_reg[1] ),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4062_ (.A1(_2270_),
    .A2(_2309_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4063_ (.A1(_1519_),
    .A2(net143),
    .B(\sense_reg[0] ),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4064_ (.A1(_2270_),
    .A2(_2310_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4065_ (.A1(_1676_),
    .A2(_2269_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4066_ (.A1(_2272_),
    .A2(net175),
    .B(\preset_n_reg[15] ),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4067_ (.A1(\state[2] ),
    .A2(_2269_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4068_ (.A1(_2312_),
    .A2(net173),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4069_ (.A1(_2278_),
    .A2(net175),
    .B(\preset_n_reg[14] ),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4070_ (.A1(net173),
    .A2(_2314_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4071_ (.A1(_2282_),
    .A2(net175),
    .B(\preset_n_reg[13] ),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4072_ (.A1(net173),
    .A2(_2315_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4073_ (.A1(_2285_),
    .A2(net175),
    .B(\preset_n_reg[12] ),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4074_ (.A1(net173),
    .A2(_2316_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4075_ (.A1(_2288_),
    .A2(net175),
    .B(\preset_n_reg[11] ),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(net173),
    .A2(_2317_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4077_ (.A1(_2291_),
    .A2(net175),
    .B(\preset_n_reg[10] ),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4078_ (.A1(net173),
    .A2(_2318_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4079_ (.A1(_2294_),
    .A2(net175),
    .B(\preset_n_reg[9] ),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(net173),
    .A2(_2319_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4081_ (.A1(_1564_),
    .A2(net176),
    .B(\preset_n_reg[8] ),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4082_ (.A1(net174),
    .A2(_2320_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4083_ (.A1(_2298_),
    .A2(net176),
    .B(\preset_n_reg[7] ),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4084_ (.A1(net174),
    .A2(_2321_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4085_ (.A1(_2301_),
    .A2(net176),
    .B(\preset_n_reg[6] ),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4086_ (.A1(net174),
    .A2(_2322_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4087_ (.A1(_2304_),
    .A2(net176),
    .B(\preset_n_reg[5] ),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4088_ (.A1(net174),
    .A2(_2323_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4089_ (.A1(_1389_),
    .A2(_2311_),
    .B(\preset_n_reg[4] ),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4090_ (.A1(_2313_),
    .A2(_2324_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4091_ (.A1(_1475_),
    .A2(_2311_),
    .B(\preset_n_reg[3] ),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(_2313_),
    .A2(_2325_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4093_ (.A1(_1533_),
    .A2(_2311_),
    .B(\preset_n_reg[2] ),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4094_ (.A1(_2313_),
    .A2(_2326_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4095_ (.A1(_1592_),
    .A2(_2311_),
    .B(\preset_n_reg[1] ),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4096_ (.A1(_2313_),
    .A2(_2327_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4097_ (.A1(_1520_),
    .A2(_2311_),
    .B(\preset_n_reg[0] ),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_2313_),
    .A2(_2328_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(net282),
    .A2(_2273_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4100_ (.A1(\col_prog_n_reg[511] ),
    .A2(net139),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4101_ (.A1(net300),
    .A2(net139),
    .B(_2330_),
    .C(net118),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4102_ (.A1(\col_prog_n_reg[510] ),
    .A2(net139),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4103_ (.A1(net298),
    .A2(net139),
    .B(_2331_),
    .C(net118),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4104_ (.A1(\col_prog_n_reg[509] ),
    .A2(net139),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4105_ (.A1(net296),
    .A2(net139),
    .B(_2332_),
    .C(net118),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4106_ (.A1(\col_prog_n_reg[508] ),
    .A2(net139),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4107_ (.A1(net293),
    .A2(net139),
    .B(_2333_),
    .C(net118),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4108_ (.A1(\col_prog_n_reg[507] ),
    .A2(net139),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4109_ (.A1(net292),
    .A2(net139),
    .B(_2334_),
    .C(net118),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4110_ (.A1(\col_prog_n_reg[506] ),
    .A2(net139),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4111_ (.A1(net290),
    .A2(net139),
    .B(_2335_),
    .C(net118),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4112_ (.A1(\col_prog_n_reg[505] ),
    .A2(net139),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4113_ (.A1(net340),
    .A2(net139),
    .B(_2336_),
    .C(net118),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4114_ (.A1(\col_prog_n_reg[504] ),
    .A2(net139),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4115_ (.A1(net338),
    .A2(net139),
    .B(_2337_),
    .C(net118),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4116_ (.A1(\col_prog_n_reg[503] ),
    .A2(net139),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4117_ (.A1(net336),
    .A2(net139),
    .B(_2338_),
    .C(net118),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4118_ (.A1(\col_prog_n_reg[502] ),
    .A2(net140),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4119_ (.A1(net334),
    .A2(net139),
    .B(_2339_),
    .C(net118),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(\col_prog_n_reg[501] ),
    .A2(net140),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4121_ (.A1(net332),
    .A2(net140),
    .B(_2340_),
    .C(net118),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4122_ (.A1(\col_prog_n_reg[500] ),
    .A2(net140),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4123_ (.A1(net329),
    .A2(net140),
    .B(_2341_),
    .C(net118),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4124_ (.A1(\col_prog_n_reg[499] ),
    .A2(net140),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4125_ (.A1(net328),
    .A2(net140),
    .B(_2342_),
    .C(net118),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4126_ (.A1(\col_prog_n_reg[498] ),
    .A2(net140),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4127_ (.A1(net326),
    .A2(net140),
    .B(_2343_),
    .C(net118),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4128_ (.A1(\col_prog_n_reg[497] ),
    .A2(net140),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4129_ (.A1(net324),
    .A2(net140),
    .B(_2344_),
    .C(net118),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4130_ (.A1(\col_prog_n_reg[496] ),
    .A2(net140),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4131_ (.A1(net321),
    .A2(net140),
    .B(_2345_),
    .C(net118),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4132_ (.A1(\col_prog_n_reg[495] ),
    .A2(net140),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4133_ (.A1(net319),
    .A2(net140),
    .B(_2346_),
    .C(net118),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4134_ (.A1(\col_prog_n_reg[494] ),
    .A2(net141),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4135_ (.A1(net317),
    .A2(net141),
    .B(_2347_),
    .C(net118),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4136_ (.A1(\col_prog_n_reg[493] ),
    .A2(net141),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4137_ (.A1(net315),
    .A2(net141),
    .B(_2348_),
    .C(net118),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(\col_prog_n_reg[492] ),
    .A2(net141),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4139_ (.A1(net313),
    .A2(net141),
    .B(_2349_),
    .C(net118),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4140_ (.A1(\col_prog_n_reg[491] ),
    .A2(net141),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4141_ (.A1(net311),
    .A2(net141),
    .B(_2350_),
    .C(net118),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(\col_prog_n_reg[490] ),
    .A2(net141),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4143_ (.A1(net309),
    .A2(net141),
    .B(_2351_),
    .C(net118),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4144_ (.A1(\col_prog_n_reg[489] ),
    .A2(net141),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4145_ (.A1(net307),
    .A2(net141),
    .B(_2352_),
    .C(net118),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4146_ (.A1(\col_prog_n_reg[488] ),
    .A2(net141),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4147_ (.A1(net304),
    .A2(net141),
    .B(_2353_),
    .C(net118),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4148_ (.A1(net282),
    .A2(\col_prog_n_reg[487] ),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4149_ (.A1(_1521_),
    .A2(_2271_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4150_ (.A1(\col_prog_n_reg[487] ),
    .A2(_2272_),
    .B1(_2355_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4151_ (.A1(_2354_),
    .A2(_2356_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4152_ (.A1(net282),
    .A2(\col_prog_n_reg[486] ),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4153_ (.A1(_1523_),
    .A2(_2271_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4154_ (.A1(\col_prog_n_reg[486] ),
    .A2(_2272_),
    .B1(_2358_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4155_ (.A1(_2357_),
    .A2(_2359_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4156_ (.A1(net282),
    .A2(\col_prog_n_reg[485] ),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4157_ (.A1(_1524_),
    .A2(_2271_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4158_ (.A1(\col_prog_n_reg[485] ),
    .A2(_2272_),
    .B1(_2361_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4159_ (.A1(_2360_),
    .A2(_2362_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4160_ (.A1(net282),
    .A2(\col_prog_n_reg[484] ),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4161_ (.A1(_1525_),
    .A2(_2271_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4162_ (.A1(\col_prog_n_reg[484] ),
    .A2(_2272_),
    .B1(_2364_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4163_ (.A1(_2363_),
    .A2(_2365_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4164_ (.A1(net282),
    .A2(\col_prog_n_reg[483] ),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4165_ (.A1(_1526_),
    .A2(_2271_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4166_ (.A1(\col_prog_n_reg[483] ),
    .A2(_2272_),
    .B1(_2367_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4167_ (.A1(_2366_),
    .A2(_2368_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4168_ (.A1(net282),
    .A2(\col_prog_n_reg[482] ),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4169_ (.A1(_1527_),
    .A2(_2271_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4170_ (.A1(\col_prog_n_reg[482] ),
    .A2(_2272_),
    .B1(_2370_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4171_ (.A1(_2369_),
    .A2(_2371_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4172_ (.A1(net282),
    .A2(\col_prog_n_reg[481] ),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4173_ (.A1(_1528_),
    .A2(_2271_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4174_ (.A1(\col_prog_n_reg[481] ),
    .A2(_2272_),
    .B1(_2373_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4175_ (.A1(_2372_),
    .A2(_2374_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4176_ (.A1(net282),
    .A2(\col_prog_n_reg[480] ),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4177_ (.A1(_1529_),
    .A2(_2271_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4178_ (.A1(\col_prog_n_reg[480] ),
    .A2(_2272_),
    .B1(_2376_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4179_ (.A1(_2375_),
    .A2(_2377_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4180_ (.A1(net282),
    .A2(net179),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(\col_prog_n_reg[479] ),
    .A2(net137),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4182_ (.A1(net300),
    .A2(net137),
    .B(_2379_),
    .C(net118),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(\col_prog_n_reg[478] ),
    .A2(net137),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4184_ (.A1(net298),
    .A2(net137),
    .B(_2380_),
    .C(net118),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4185_ (.A1(\col_prog_n_reg[477] ),
    .A2(net137),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4186_ (.A1(net296),
    .A2(net137),
    .B(_2381_),
    .C(net118),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(\col_prog_n_reg[476] ),
    .A2(net137),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4188_ (.A1(net293),
    .A2(net137),
    .B(_2382_),
    .C(net118),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(\col_prog_n_reg[475] ),
    .A2(net137),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4190_ (.A1(net292),
    .A2(net137),
    .B(_2383_),
    .C(net118),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(\col_prog_n_reg[474] ),
    .A2(net137),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4192_ (.A1(net290),
    .A2(net137),
    .B(_2384_),
    .C(net118),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4193_ (.A1(\col_prog_n_reg[473] ),
    .A2(net137),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4194_ (.A1(net340),
    .A2(net137),
    .B(_2385_),
    .C(net118),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4195_ (.A1(\col_prog_n_reg[472] ),
    .A2(net137),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4196_ (.A1(net338),
    .A2(net137),
    .B(_2386_),
    .C(net118),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(\col_prog_n_reg[471] ),
    .A2(net137),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4198_ (.A1(net336),
    .A2(net137),
    .B(_2387_),
    .C(net118),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4199_ (.A1(\col_prog_n_reg[470] ),
    .A2(net137),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4200_ (.A1(net334),
    .A2(net137),
    .B(_2388_),
    .C(net118),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4201_ (.A1(\col_prog_n_reg[469] ),
    .A2(net138),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4202_ (.A1(net332),
    .A2(net138),
    .B(_2389_),
    .C(net118),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4203_ (.A1(\col_prog_n_reg[468] ),
    .A2(net138),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4204_ (.A1(net329),
    .A2(net138),
    .B(_2390_),
    .C(net118),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4205_ (.A1(\col_prog_n_reg[467] ),
    .A2(net138),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4206_ (.A1(net328),
    .A2(net138),
    .B(_2391_),
    .C(net118),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4207_ (.A1(\col_prog_n_reg[466] ),
    .A2(net138),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4208_ (.A1(net326),
    .A2(net138),
    .B(_2392_),
    .C(net118),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(\col_prog_n_reg[465] ),
    .A2(net138),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4210_ (.A1(net324),
    .A2(net138),
    .B(_2393_),
    .C(net118),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4211_ (.A1(\col_prog_n_reg[464] ),
    .A2(net138),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4212_ (.A1(net321),
    .A2(net138),
    .B(_2394_),
    .C(net118),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4213_ (.A1(\col_prog_n_reg[463] ),
    .A2(net138),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4214_ (.A1(net319),
    .A2(net138),
    .B(_2395_),
    .C(net118),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4215_ (.A1(\col_prog_n_reg[462] ),
    .A2(net138),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4216_ (.A1(net317),
    .A2(net138),
    .B(_2396_),
    .C(net118),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4217_ (.A1(\col_prog_n_reg[461] ),
    .A2(_2378_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4218_ (.A1(net315),
    .A2(_2378_),
    .B(_2397_),
    .C(net118),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4219_ (.A1(\col_prog_n_reg[460] ),
    .A2(_2378_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4220_ (.A1(net313),
    .A2(_2378_),
    .B(_2398_),
    .C(net118),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4221_ (.A1(\col_prog_n_reg[459] ),
    .A2(_2378_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4222_ (.A1(net311),
    .A2(_2378_),
    .B(_2399_),
    .C(net118),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4223_ (.A1(\col_prog_n_reg[458] ),
    .A2(_2378_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4224_ (.A1(net309),
    .A2(_2378_),
    .B(_2400_),
    .C(net118),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4225_ (.A1(\col_prog_n_reg[457] ),
    .A2(_2378_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4226_ (.A1(net307),
    .A2(_2378_),
    .B(_2401_),
    .C(net118),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4227_ (.A1(\col_prog_n_reg[456] ),
    .A2(_2378_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4228_ (.A1(net304),
    .A2(_2378_),
    .B(_2402_),
    .C(net118),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4229_ (.A1(net282),
    .A2(\col_prog_n_reg[455] ),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4230_ (.A1(_1521_),
    .A2(_2276_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4231_ (.A1(\col_prog_n_reg[455] ),
    .A2(_2278_),
    .B1(_2404_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4232_ (.A1(_2403_),
    .A2(_2405_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4233_ (.A1(net282),
    .A2(\col_prog_n_reg[454] ),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4234_ (.A1(_1523_),
    .A2(_2276_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4235_ (.A1(\col_prog_n_reg[454] ),
    .A2(_2278_),
    .B1(_2407_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4236_ (.A1(_2406_),
    .A2(_2408_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4237_ (.A1(net282),
    .A2(\col_prog_n_reg[453] ),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4238_ (.A1(_1524_),
    .A2(_2276_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4239_ (.A1(\col_prog_n_reg[453] ),
    .A2(_2278_),
    .B1(_2410_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4240_ (.A1(_2409_),
    .A2(_2411_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4241_ (.A1(net282),
    .A2(\col_prog_n_reg[452] ),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4242_ (.A1(_1525_),
    .A2(_2276_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4243_ (.A1(\col_prog_n_reg[452] ),
    .A2(_2278_),
    .B1(_2413_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4244_ (.A1(_2412_),
    .A2(_2414_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4245_ (.A1(net282),
    .A2(\col_prog_n_reg[451] ),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4246_ (.A1(_1526_),
    .A2(_2276_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4247_ (.A1(\col_prog_n_reg[451] ),
    .A2(_2278_),
    .B1(_2416_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4248_ (.A1(_2415_),
    .A2(_2417_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4249_ (.A1(net282),
    .A2(\col_prog_n_reg[450] ),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4250_ (.A1(_1527_),
    .A2(_2276_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4251_ (.A1(\col_prog_n_reg[450] ),
    .A2(_2278_),
    .B1(_2419_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4252_ (.A1(_2418_),
    .A2(_2420_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4253_ (.A1(net282),
    .A2(\col_prog_n_reg[449] ),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4254_ (.A1(_1528_),
    .A2(_2276_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4255_ (.A1(\col_prog_n_reg[449] ),
    .A2(_2278_),
    .B1(_2422_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4256_ (.A1(_2421_),
    .A2(_2423_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4257_ (.A1(net282),
    .A2(\col_prog_n_reg[448] ),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4258_ (.A1(_1529_),
    .A2(_2276_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4259_ (.A1(\col_prog_n_reg[448] ),
    .A2(_2278_),
    .B1(_2425_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4260_ (.A1(_2424_),
    .A2(_2426_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4261_ (.A1(net282),
    .A2(net178),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4262_ (.A1(\col_prog_n_reg[447] ),
    .A2(net135),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4263_ (.A1(net300),
    .A2(net135),
    .B(_2428_),
    .C(net118),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4264_ (.A1(\col_prog_n_reg[446] ),
    .A2(net135),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4265_ (.A1(net298),
    .A2(net135),
    .B(_2429_),
    .C(net118),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4266_ (.A1(\col_prog_n_reg[445] ),
    .A2(net135),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4267_ (.A1(net296),
    .A2(net135),
    .B(_2430_),
    .C(net118),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4268_ (.A1(\col_prog_n_reg[444] ),
    .A2(net135),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4269_ (.A1(net293),
    .A2(net135),
    .B(_2431_),
    .C(net118),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4270_ (.A1(\col_prog_n_reg[443] ),
    .A2(net135),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4271_ (.A1(net292),
    .A2(net135),
    .B(_2432_),
    .C(net118),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4272_ (.A1(\col_prog_n_reg[442] ),
    .A2(net135),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4273_ (.A1(net290),
    .A2(net135),
    .B(_2433_),
    .C(net118),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4274_ (.A1(\col_prog_n_reg[441] ),
    .A2(net135),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4275_ (.A1(net340),
    .A2(net135),
    .B(_2434_),
    .C(net118),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4276_ (.A1(\col_prog_n_reg[440] ),
    .A2(net135),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4277_ (.A1(net338),
    .A2(net135),
    .B(_2435_),
    .C(net118),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4278_ (.A1(\col_prog_n_reg[439] ),
    .A2(net135),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4279_ (.A1(net336),
    .A2(net135),
    .B(_2436_),
    .C(net118),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4280_ (.A1(\col_prog_n_reg[438] ),
    .A2(net135),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4281_ (.A1(net334),
    .A2(net135),
    .B(_2437_),
    .C(net118),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(\col_prog_n_reg[437] ),
    .A2(net136),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4283_ (.A1(net332),
    .A2(net136),
    .B(_2438_),
    .C(net118),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4284_ (.A1(\col_prog_n_reg[436] ),
    .A2(net136),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4285_ (.A1(net329),
    .A2(net136),
    .B(_2439_),
    .C(net118),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4286_ (.A1(\col_prog_n_reg[435] ),
    .A2(net136),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4287_ (.A1(net328),
    .A2(net136),
    .B(_2440_),
    .C(net118),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4288_ (.A1(\col_prog_n_reg[434] ),
    .A2(net136),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4289_ (.A1(net326),
    .A2(net136),
    .B(_2441_),
    .C(net118),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4290_ (.A1(\col_prog_n_reg[433] ),
    .A2(net136),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4291_ (.A1(net324),
    .A2(net136),
    .B(_2442_),
    .C(net118),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(\col_prog_n_reg[432] ),
    .A2(net136),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4293_ (.A1(net321),
    .A2(net136),
    .B(_2443_),
    .C(net118),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4294_ (.A1(\col_prog_n_reg[431] ),
    .A2(net136),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4295_ (.A1(net319),
    .A2(net136),
    .B(_2444_),
    .C(net118),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(\col_prog_n_reg[430] ),
    .A2(_2427_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4297_ (.A1(net317),
    .A2(_2427_),
    .B(_2445_),
    .C(net118),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4298_ (.A1(\col_prog_n_reg[429] ),
    .A2(_2427_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4299_ (.A1(net315),
    .A2(_2427_),
    .B(_2446_),
    .C(net118),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4300_ (.A1(\col_prog_n_reg[428] ),
    .A2(_2427_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4301_ (.A1(net313),
    .A2(_2427_),
    .B(_2447_),
    .C(net118),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4302_ (.A1(\col_prog_n_reg[427] ),
    .A2(_2427_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4303_ (.A1(net311),
    .A2(_2427_),
    .B(_2448_),
    .C(net118),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4304_ (.A1(\col_prog_n_reg[426] ),
    .A2(_2427_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4305_ (.A1(net309),
    .A2(_2427_),
    .B(_2449_),
    .C(net118),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4306_ (.A1(\col_prog_n_reg[425] ),
    .A2(_2427_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4307_ (.A1(net307),
    .A2(_2427_),
    .B(_2450_),
    .C(net118),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(\col_prog_n_reg[424] ),
    .A2(_2427_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4309_ (.A1(net304),
    .A2(_2427_),
    .B(_2451_),
    .C(net118),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4310_ (.A1(net282),
    .A2(\col_prog_n_reg[423] ),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4311_ (.A1(_1521_),
    .A2(net257),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4312_ (.A1(\col_prog_n_reg[423] ),
    .A2(_2282_),
    .B1(net134),
    .B2(_1566_),
    .C(net164),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4313_ (.A1(_2452_),
    .A2(_2454_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4314_ (.A1(net282),
    .A2(\col_prog_n_reg[422] ),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4315_ (.A1(_1523_),
    .A2(net257),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4316_ (.A1(\col_prog_n_reg[422] ),
    .A2(_2282_),
    .B1(_2456_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4317_ (.A1(_2455_),
    .A2(_2457_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4318_ (.A1(net282),
    .A2(\col_prog_n_reg[421] ),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4319_ (.A1(_1524_),
    .A2(net257),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4320_ (.A1(\col_prog_n_reg[421] ),
    .A2(_2282_),
    .B1(_2459_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4321_ (.A1(_2458_),
    .A2(_2460_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4322_ (.A1(net282),
    .A2(\col_prog_n_reg[420] ),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4323_ (.A1(_1525_),
    .A2(net257),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4324_ (.A1(\col_prog_n_reg[420] ),
    .A2(_2282_),
    .B1(_2462_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4325_ (.A1(_2461_),
    .A2(_2463_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4326_ (.A1(net282),
    .A2(\col_prog_n_reg[419] ),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4327_ (.A1(_1526_),
    .A2(net257),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4328_ (.A1(\col_prog_n_reg[419] ),
    .A2(_2282_),
    .B1(_2465_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(_2464_),
    .A2(_2466_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4330_ (.A1(net282),
    .A2(\col_prog_n_reg[418] ),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4331_ (.A1(_1527_),
    .A2(net257),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4332_ (.A1(\col_prog_n_reg[418] ),
    .A2(_2282_),
    .B1(_2468_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4333_ (.A1(_2467_),
    .A2(_2469_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4334_ (.A1(net282),
    .A2(\col_prog_n_reg[417] ),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4335_ (.A1(_1528_),
    .A2(net257),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4336_ (.A1(\col_prog_n_reg[417] ),
    .A2(_2282_),
    .B1(_2471_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4337_ (.A1(_2470_),
    .A2(_2472_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4338_ (.A1(net282),
    .A2(\col_prog_n_reg[416] ),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4339_ (.A1(_1529_),
    .A2(net257),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4340_ (.A1(\col_prog_n_reg[416] ),
    .A2(_2282_),
    .B1(_2474_),
    .B2(_1566_),
    .C(net164),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4341_ (.A1(_2473_),
    .A2(_2475_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4342_ (.A1(_1309_),
    .A2(_2285_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4343_ (.A1(net282),
    .A2(_2284_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(net300),
    .A2(net170),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4345_ (.A1(\col_prog_n_reg[415] ),
    .A2(net170),
    .B(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4346_ (.A1(net119),
    .A2(_2479_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4347_ (.A1(net298),
    .A2(net170),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4348_ (.A1(\col_prog_n_reg[414] ),
    .A2(net170),
    .B(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4349_ (.A1(net119),
    .A2(_2481_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4350_ (.A1(net296),
    .A2(net170),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4351_ (.A1(\col_prog_n_reg[413] ),
    .A2(net170),
    .B(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(net119),
    .A2(_2483_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4353_ (.A1(net293),
    .A2(net170),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4354_ (.A1(\col_prog_n_reg[412] ),
    .A2(net170),
    .B(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4355_ (.A1(net119),
    .A2(_2485_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4356_ (.A1(net292),
    .A2(net170),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4357_ (.A1(\col_prog_n_reg[411] ),
    .A2(net170),
    .B(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4358_ (.A1(net119),
    .A2(_2487_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4359_ (.A1(net290),
    .A2(net170),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4360_ (.A1(\col_prog_n_reg[410] ),
    .A2(net170),
    .B(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4361_ (.A1(net119),
    .A2(_2489_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4362_ (.A1(\col_prog_n_reg[409] ),
    .A2(net133),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4363_ (.A1(net340),
    .A2(net133),
    .B(_2490_),
    .C(net119),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4364_ (.A1(\col_prog_n_reg[408] ),
    .A2(net133),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4365_ (.A1(net338),
    .A2(net133),
    .B(_2491_),
    .C(net119),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4366_ (.A1(\col_prog_n_reg[407] ),
    .A2(net133),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4367_ (.A1(net336),
    .A2(net133),
    .B(_2492_),
    .C(net119),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(\col_prog_n_reg[406] ),
    .A2(net133),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4369_ (.A1(net334),
    .A2(net133),
    .B(_2493_),
    .C(net119),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4370_ (.A1(\col_prog_n_reg[405] ),
    .A2(net133),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4371_ (.A1(net332),
    .A2(net133),
    .B(_2494_),
    .C(net119),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(\col_prog_n_reg[404] ),
    .A2(net133),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4373_ (.A1(net329),
    .A2(net133),
    .B(_2495_),
    .C(net119),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4374_ (.A1(\col_prog_n_reg[403] ),
    .A2(net133),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4375_ (.A1(net328),
    .A2(net133),
    .B(_2496_),
    .C(net119),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4376_ (.A1(\col_prog_n_reg[402] ),
    .A2(net133),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4377_ (.A1(net326),
    .A2(net133),
    .B(_2497_),
    .C(net119),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(\col_prog_n_reg[401] ),
    .A2(net133),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4379_ (.A1(net324),
    .A2(net133),
    .B(_2498_),
    .C(net119),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4380_ (.A1(\col_prog_n_reg[400] ),
    .A2(net133),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4381_ (.A1(net321),
    .A2(net133),
    .B(_2499_),
    .C(net119),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4382_ (.A1(\col_prog_n_reg[399] ),
    .A2(_2477_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4383_ (.A1(net319),
    .A2(_2477_),
    .B(_2500_),
    .C(net119),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4384_ (.A1(\col_prog_n_reg[398] ),
    .A2(_2477_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4385_ (.A1(net317),
    .A2(_2477_),
    .B(_2501_),
    .C(net119),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(\col_prog_n_reg[397] ),
    .A2(_2477_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4387_ (.A1(net315),
    .A2(_2477_),
    .B(_2502_),
    .C(net119),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4388_ (.A1(\col_prog_n_reg[396] ),
    .A2(_2477_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4389_ (.A1(net313),
    .A2(_2477_),
    .B(_2503_),
    .C(net119),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(\col_prog_n_reg[395] ),
    .A2(_2477_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4391_ (.A1(net311),
    .A2(_2477_),
    .B(_2504_),
    .C(net119),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4392_ (.A1(\col_prog_n_reg[394] ),
    .A2(_2477_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4393_ (.A1(net309),
    .A2(_2477_),
    .B(_2505_),
    .C(net119),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4394_ (.A1(\col_prog_n_reg[393] ),
    .A2(_2477_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4395_ (.A1(net307),
    .A2(_2477_),
    .B(_2506_),
    .C(net118),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(\col_prog_n_reg[392] ),
    .A2(_2477_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4397_ (.A1(net304),
    .A2(_2477_),
    .B(_2507_),
    .C(net118),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4398_ (.A1(net167),
    .A2(net172),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4399_ (.A1(\col_prog_n_reg[391] ),
    .A2(net167),
    .A3(net172),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4400_ (.A1(\col_prog_n_reg[391] ),
    .A2(_2285_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4401_ (.A1(net115),
    .A2(_2509_),
    .B(_2510_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4402_ (.A1(net113),
    .A2(net172),
    .B1(_2508_),
    .B2(_1349_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4403_ (.A1(net111),
    .A2(net172),
    .B1(_2508_),
    .B2(_1350_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4404_ (.A1(net109),
    .A2(net172),
    .B1(_2508_),
    .B2(_1351_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4405_ (.A1(net107),
    .A2(net172),
    .B1(_2508_),
    .B2(_1352_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4406_ (.A1(net105),
    .A2(net177),
    .B1(_2508_),
    .B2(_1353_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4407_ (.A1(net103),
    .A2(net172),
    .B1(_2508_),
    .B2(_1354_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4408_ (.A1(net101),
    .A2(net172),
    .B1(_2508_),
    .B2(_1355_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4409_ (.A1(_1309_),
    .A2(_2288_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4410_ (.A1(net282),
    .A2(net256),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4411_ (.A1(\col_prog_n_reg[383] ),
    .A2(net168),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4412_ (.A1(net300),
    .A2(net168),
    .B(_2513_),
    .C(net119),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(\col_prog_n_reg[382] ),
    .A2(net168),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4414_ (.A1(net298),
    .A2(net168),
    .B(_2514_),
    .C(net119),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4415_ (.A1(\col_prog_n_reg[381] ),
    .A2(net168),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4416_ (.A1(net296),
    .A2(net168),
    .B(_2515_),
    .C(net119),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(\col_prog_n_reg[380] ),
    .A2(net168),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4418_ (.A1(net293),
    .A2(net168),
    .B(_2516_),
    .C(net119),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(\col_prog_n_reg[379] ),
    .A2(net168),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4420_ (.A1(net292),
    .A2(net168),
    .B(_2517_),
    .C(net119),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4421_ (.A1(\col_prog_n_reg[378] ),
    .A2(net168),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4422_ (.A1(net290),
    .A2(net168),
    .B(_2518_),
    .C(net119),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(\col_prog_n_reg[377] ),
    .A2(net168),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4424_ (.A1(net340),
    .A2(net168),
    .B(_2519_),
    .C(net119),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4425_ (.A1(\col_prog_n_reg[376] ),
    .A2(net168),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4426_ (.A1(net338),
    .A2(net168),
    .B(_2520_),
    .C(net119),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4427_ (.A1(\col_prog_n_reg[375] ),
    .A2(net168),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4428_ (.A1(net336),
    .A2(net168),
    .B(_2521_),
    .C(net119),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4429_ (.A1(\col_prog_n_reg[374] ),
    .A2(net168),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4430_ (.A1(net334),
    .A2(net168),
    .B(_2522_),
    .C(net119),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4431_ (.A1(\col_prog_n_reg[373] ),
    .A2(net169),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4432_ (.A1(net332),
    .A2(net168),
    .B(_2523_),
    .C(net119),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(\col_prog_n_reg[372] ),
    .A2(net169),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4434_ (.A1(net329),
    .A2(net169),
    .B(_2524_),
    .C(net119),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4435_ (.A1(\col_prog_n_reg[371] ),
    .A2(net169),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4436_ (.A1(net328),
    .A2(net169),
    .B(_2525_),
    .C(net119),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(\col_prog_n_reg[370] ),
    .A2(net169),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4438_ (.A1(net326),
    .A2(net169),
    .B(_2526_),
    .C(net119),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(\col_prog_n_reg[369] ),
    .A2(net169),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4440_ (.A1(net324),
    .A2(net169),
    .B(_2527_),
    .C(net119),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(\col_prog_n_reg[368] ),
    .A2(net169),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4442_ (.A1(net321),
    .A2(net169),
    .B(_2528_),
    .C(net119),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4443_ (.A1(\col_prog_n_reg[367] ),
    .A2(net169),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4444_ (.A1(net319),
    .A2(net169),
    .B(_2529_),
    .C(net119),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4445_ (.A1(\col_prog_n_reg[366] ),
    .A2(net169),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4446_ (.A1(net317),
    .A2(net169),
    .B(_2530_),
    .C(net119),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4447_ (.A1(\col_prog_n_reg[365] ),
    .A2(net169),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4448_ (.A1(net315),
    .A2(net169),
    .B(_2531_),
    .C(net119),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4449_ (.A1(\col_prog_n_reg[364] ),
    .A2(_2512_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4450_ (.A1(net313),
    .A2(_2512_),
    .B(_2532_),
    .C(net119),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4451_ (.A1(\col_prog_n_reg[363] ),
    .A2(_2512_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4452_ (.A1(net311),
    .A2(_2512_),
    .B(_2533_),
    .C(net119),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(\col_prog_n_reg[362] ),
    .A2(_2512_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4454_ (.A1(net309),
    .A2(_2512_),
    .B(_2534_),
    .C(net119),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(\col_prog_n_reg[361] ),
    .A2(_2512_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4456_ (.A1(net307),
    .A2(_2512_),
    .B(_2535_),
    .C(net119),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4457_ (.A1(\col_prog_n_reg[360] ),
    .A2(_2512_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4458_ (.A1(net304),
    .A2(_2512_),
    .B(_2536_),
    .C(net119),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4459_ (.A1(net167),
    .A2(_2511_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4460_ (.A1(\col_prog_n_reg[359] ),
    .A2(net167),
    .A3(_2511_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4461_ (.A1(\col_prog_n_reg[359] ),
    .A2(_2288_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4462_ (.A1(net115),
    .A2(_2538_),
    .B(_2539_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4463_ (.A1(net113),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1356_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4464_ (.A1(net111),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1357_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4465_ (.A1(net109),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1358_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4466_ (.A1(net107),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1359_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4467_ (.A1(net105),
    .A2(net255),
    .B1(_2537_),
    .B2(_1360_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4468_ (.A1(net103),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1361_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4469_ (.A1(net101),
    .A2(_2511_),
    .B1(_2537_),
    .B2(_1362_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4470_ (.A1(net282),
    .A2(_2290_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4471_ (.A1(\col_prog_n_reg[351] ),
    .A2(net131),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4472_ (.A1(net300),
    .A2(net131),
    .B(_2541_),
    .C(net120),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4473_ (.A1(\col_prog_n_reg[350] ),
    .A2(net131),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4474_ (.A1(net298),
    .A2(net131),
    .B(_2542_),
    .C(net120),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4475_ (.A1(\col_prog_n_reg[349] ),
    .A2(net131),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4476_ (.A1(net296),
    .A2(net131),
    .B(_2543_),
    .C(net120),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4477_ (.A1(\col_prog_n_reg[348] ),
    .A2(net131),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4478_ (.A1(net293),
    .A2(net131),
    .B(_2544_),
    .C(net120),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4479_ (.A1(\col_prog_n_reg[347] ),
    .A2(net131),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4480_ (.A1(net292),
    .A2(net131),
    .B(_2545_),
    .C(net120),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4481_ (.A1(\col_prog_n_reg[346] ),
    .A2(net131),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4482_ (.A1(net290),
    .A2(net131),
    .B(_2546_),
    .C(net120),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4483_ (.A1(\col_prog_n_reg[345] ),
    .A2(net131),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4484_ (.A1(net340),
    .A2(net131),
    .B(_2547_),
    .C(net120),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(\col_prog_n_reg[344] ),
    .A2(net131),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4486_ (.A1(net338),
    .A2(net131),
    .B(_2548_),
    .C(net120),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4487_ (.A1(\col_prog_n_reg[343] ),
    .A2(net131),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4488_ (.A1(net336),
    .A2(net131),
    .B(_2549_),
    .C(net120),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4489_ (.A1(\col_prog_n_reg[342] ),
    .A2(net131),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4490_ (.A1(net334),
    .A2(net131),
    .B(_2550_),
    .C(net120),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4491_ (.A1(\col_prog_n_reg[341] ),
    .A2(net132),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4492_ (.A1(net332),
    .A2(net132),
    .B(_2551_),
    .C(net120),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(\col_prog_n_reg[340] ),
    .A2(net132),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4494_ (.A1(net329),
    .A2(net132),
    .B(_2552_),
    .C(net120),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4495_ (.A1(\col_prog_n_reg[339] ),
    .A2(net132),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4496_ (.A1(net328),
    .A2(net132),
    .B(_2553_),
    .C(net120),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4497_ (.A1(\col_prog_n_reg[338] ),
    .A2(net132),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4498_ (.A1(net326),
    .A2(net132),
    .B(_2554_),
    .C(net120),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4499_ (.A1(\col_prog_n_reg[337] ),
    .A2(net132),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4500_ (.A1(net324),
    .A2(net132),
    .B(_2555_),
    .C(net120),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4501_ (.A1(\col_prog_n_reg[336] ),
    .A2(net132),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4502_ (.A1(net321),
    .A2(net132),
    .B(_2556_),
    .C(net120),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(\col_prog_n_reg[335] ),
    .A2(net132),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4504_ (.A1(net319),
    .A2(net132),
    .B(_2557_),
    .C(net120),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4505_ (.A1(\col_prog_n_reg[334] ),
    .A2(_2540_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4506_ (.A1(net317),
    .A2(_2540_),
    .B(_2558_),
    .C(net120),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4507_ (.A1(\col_prog_n_reg[333] ),
    .A2(_2540_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4508_ (.A1(net315),
    .A2(_2540_),
    .B(_2559_),
    .C(net120),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4509_ (.A1(\col_prog_n_reg[332] ),
    .A2(_2540_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4510_ (.A1(net313),
    .A2(_2540_),
    .B(_2560_),
    .C(net120),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4511_ (.A1(\col_prog_n_reg[331] ),
    .A2(_2540_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4512_ (.A1(net311),
    .A2(_2540_),
    .B(_2561_),
    .C(net120),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4513_ (.A1(\col_prog_n_reg[330] ),
    .A2(_2540_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4514_ (.A1(net309),
    .A2(_2540_),
    .B(_2562_),
    .C(net120),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4515_ (.A1(\col_prog_n_reg[329] ),
    .A2(_2540_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4516_ (.A1(net307),
    .A2(_2540_),
    .B(_2563_),
    .C(net119),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4517_ (.A1(\col_prog_n_reg[328] ),
    .A2(_2540_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4518_ (.A1(net304),
    .A2(_2540_),
    .B(_2564_),
    .C(net119),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4519_ (.A1(net282),
    .A2(\col_prog_n_reg[327] ),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4520_ (.A1(_1563_),
    .A2(_1566_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[327] ),
    .C(net165),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4521_ (.A1(_2565_),
    .A2(_2566_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4522_ (.A1(net282),
    .A2(\col_prog_n_reg[326] ),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4523_ (.A1(_1566_),
    .A2(_1569_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[326] ),
    .C(net165),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4524_ (.A1(_2567_),
    .A2(_2568_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4525_ (.A1(net282),
    .A2(\col_prog_n_reg[325] ),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4526_ (.A1(_1566_),
    .A2(_1572_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[325] ),
    .C(net165),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4527_ (.A1(_2569_),
    .A2(_2570_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4528_ (.A1(net282),
    .A2(\col_prog_n_reg[324] ),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4529_ (.A1(_1566_),
    .A2(_1575_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[324] ),
    .C(net165),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4530_ (.A1(_2571_),
    .A2(_2572_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4531_ (.A1(net282),
    .A2(\col_prog_n_reg[323] ),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4532_ (.A1(_1566_),
    .A2(_1578_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[323] ),
    .C(net165),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4533_ (.A1(_2573_),
    .A2(_2574_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4534_ (.A1(net282),
    .A2(\col_prog_n_reg[322] ),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4535_ (.A1(_1566_),
    .A2(_1581_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[322] ),
    .C(net165),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4536_ (.A1(_2575_),
    .A2(_2576_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4537_ (.A1(net282),
    .A2(\col_prog_n_reg[321] ),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4538_ (.A1(_1566_),
    .A2(_1584_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[321] ),
    .C(net165),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4539_ (.A1(_2577_),
    .A2(_2578_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4540_ (.A1(net282),
    .A2(\col_prog_n_reg[320] ),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4541_ (.A1(_1566_),
    .A2(_1587_),
    .B1(_2291_),
    .B2(\col_prog_n_reg[320] ),
    .C(net165),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4542_ (.A1(_2579_),
    .A2(_2580_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4543_ (.A1(net282),
    .A2(_2293_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4544_ (.A1(\col_prog_n_reg[319] ),
    .A2(net129),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4545_ (.A1(net300),
    .A2(net129),
    .B(_2582_),
    .C(net120),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4546_ (.A1(\col_prog_n_reg[318] ),
    .A2(net129),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4547_ (.A1(net298),
    .A2(net129),
    .B(_2583_),
    .C(net120),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4548_ (.A1(\col_prog_n_reg[317] ),
    .A2(net129),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4549_ (.A1(net296),
    .A2(net129),
    .B(_2584_),
    .C(net120),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4550_ (.A1(\col_prog_n_reg[316] ),
    .A2(net129),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4551_ (.A1(net293),
    .A2(net129),
    .B(_2585_),
    .C(net120),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4552_ (.A1(\col_prog_n_reg[315] ),
    .A2(net129),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4553_ (.A1(net292),
    .A2(net129),
    .B(_2586_),
    .C(net120),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4554_ (.A1(\col_prog_n_reg[314] ),
    .A2(net129),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4555_ (.A1(net290),
    .A2(net129),
    .B(_2587_),
    .C(net120),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4556_ (.A1(\col_prog_n_reg[313] ),
    .A2(net129),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4557_ (.A1(net340),
    .A2(net129),
    .B(_2588_),
    .C(net120),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4558_ (.A1(\col_prog_n_reg[312] ),
    .A2(net129),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4559_ (.A1(net338),
    .A2(net129),
    .B(_2589_),
    .C(net120),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4560_ (.A1(\col_prog_n_reg[311] ),
    .A2(net129),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4561_ (.A1(net336),
    .A2(net129),
    .B(_2590_),
    .C(net120),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4562_ (.A1(\col_prog_n_reg[310] ),
    .A2(net129),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4563_ (.A1(net334),
    .A2(net129),
    .B(_2591_),
    .C(net120),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(\col_prog_n_reg[309] ),
    .A2(net130),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4565_ (.A1(net332),
    .A2(net129),
    .B(_2592_),
    .C(net120),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4566_ (.A1(\col_prog_n_reg[308] ),
    .A2(net130),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4567_ (.A1(net329),
    .A2(net130),
    .B(_2593_),
    .C(net120),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4568_ (.A1(\col_prog_n_reg[307] ),
    .A2(net130),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4569_ (.A1(net328),
    .A2(net130),
    .B(_2594_),
    .C(net120),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4570_ (.A1(\col_prog_n_reg[306] ),
    .A2(net130),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4571_ (.A1(net326),
    .A2(net130),
    .B(_2595_),
    .C(net120),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(\col_prog_n_reg[305] ),
    .A2(net130),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4573_ (.A1(net324),
    .A2(net130),
    .B(_2596_),
    .C(net120),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4574_ (.A1(\col_prog_n_reg[304] ),
    .A2(net130),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4575_ (.A1(net321),
    .A2(net130),
    .B(_2597_),
    .C(net120),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(\col_prog_n_reg[303] ),
    .A2(net130),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4577_ (.A1(net319),
    .A2(net130),
    .B(_2598_),
    .C(net120),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4578_ (.A1(\col_prog_n_reg[302] ),
    .A2(net130),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4579_ (.A1(net317),
    .A2(net130),
    .B(_2599_),
    .C(net120),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4580_ (.A1(\col_prog_n_reg[301] ),
    .A2(_2581_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4581_ (.A1(net315),
    .A2(_2581_),
    .B(_2600_),
    .C(net120),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(\col_prog_n_reg[300] ),
    .A2(_2581_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4583_ (.A1(net313),
    .A2(_2581_),
    .B(_2601_),
    .C(net120),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(\col_prog_n_reg[299] ),
    .A2(_2581_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4585_ (.A1(net311),
    .A2(_2581_),
    .B(_2602_),
    .C(net120),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4586_ (.A1(\col_prog_n_reg[298] ),
    .A2(_2581_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4587_ (.A1(net309),
    .A2(_2581_),
    .B(_2603_),
    .C(net120),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(\col_prog_n_reg[297] ),
    .A2(_2581_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4589_ (.A1(net307),
    .A2(_2581_),
    .B(_2604_),
    .C(net120),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(\col_prog_n_reg[296] ),
    .A2(_2581_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4591_ (.A1(net304),
    .A2(_2581_),
    .B(_2605_),
    .C(net120),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4592_ (.A1(net282),
    .A2(\col_prog_n_reg[295] ),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4593_ (.A1(_1566_),
    .A2(_1619_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[295] ),
    .C(net165),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4594_ (.A1(_2606_),
    .A2(_2607_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4595_ (.A1(net282),
    .A2(\col_prog_n_reg[294] ),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4596_ (.A1(_1566_),
    .A2(_1622_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[294] ),
    .C(net165),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4597_ (.A1(_2608_),
    .A2(_2609_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4598_ (.A1(net282),
    .A2(\col_prog_n_reg[293] ),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4599_ (.A1(_1566_),
    .A2(_1625_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[293] ),
    .C(net165),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4600_ (.A1(_2610_),
    .A2(_2611_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4601_ (.A1(net282),
    .A2(\col_prog_n_reg[292] ),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4602_ (.A1(_1566_),
    .A2(_1628_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[292] ),
    .C(net165),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4603_ (.A1(_2612_),
    .A2(_2613_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4604_ (.A1(net282),
    .A2(\col_prog_n_reg[291] ),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4605_ (.A1(_1566_),
    .A2(_1631_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[291] ),
    .C(net165),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4606_ (.A1(_2614_),
    .A2(_2615_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4607_ (.A1(net282),
    .A2(\col_prog_n_reg[290] ),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4608_ (.A1(_1566_),
    .A2(_1634_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[290] ),
    .C(net165),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4609_ (.A1(_2616_),
    .A2(_2617_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4610_ (.A1(net282),
    .A2(\col_prog_n_reg[289] ),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4611_ (.A1(_1566_),
    .A2(_1637_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[289] ),
    .C(net165),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4612_ (.A1(_2618_),
    .A2(_2619_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4613_ (.A1(net282),
    .A2(\col_prog_n_reg[288] ),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4614_ (.A1(_1566_),
    .A2(_1640_),
    .B1(_2294_),
    .B2(\col_prog_n_reg[288] ),
    .C(net165),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4615_ (.A1(_2620_),
    .A2(_2621_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4616_ (.A1(\state[3] ),
    .A2(net360),
    .A3(net287),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4617_ (.A1(\col_prog_n_reg[287] ),
    .A2(net253),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4618_ (.A1(_1478_),
    .A2(net253),
    .B(_2623_),
    .C(net121),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(\col_prog_n_reg[286] ),
    .A2(net253),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4620_ (.A1(_1481_),
    .A2(net253),
    .B(_2624_),
    .C(net121),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(\col_prog_n_reg[285] ),
    .A2(net253),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4622_ (.A1(_1484_),
    .A2(net253),
    .B(_2625_),
    .C(net121),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4623_ (.A1(\col_prog_n_reg[284] ),
    .A2(net253),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4624_ (.A1(_1487_),
    .A2(net253),
    .B(_2626_),
    .C(net121),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4625_ (.A1(\col_prog_n_reg[283] ),
    .A2(net253),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4626_ (.A1(_1490_),
    .A2(net253),
    .B(_2627_),
    .C(net121),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(\col_prog_n_reg[282] ),
    .A2(net253),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4628_ (.A1(_1493_),
    .A2(net253),
    .B(_2628_),
    .C(net121),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4629_ (.A1(\col_prog_n_reg[281] ),
    .A2(net253),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4630_ (.A1(_1392_),
    .A2(net253),
    .B(_2629_),
    .C(net121),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(\col_prog_n_reg[280] ),
    .A2(net253),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4632_ (.A1(_1395_),
    .A2(net253),
    .B(_2630_),
    .C(net121),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4633_ (.A1(\col_prog_n_reg[279] ),
    .A2(net253),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4634_ (.A1(_1398_),
    .A2(net253),
    .B(_2631_),
    .C(net121),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(\col_prog_n_reg[278] ),
    .A2(net253),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4636_ (.A1(_1401_),
    .A2(net253),
    .B(_2632_),
    .C(net121),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4637_ (.A1(\col_prog_n_reg[277] ),
    .A2(net253),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4638_ (.A1(_1404_),
    .A2(net253),
    .B(_2633_),
    .C(net121),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(\col_prog_n_reg[276] ),
    .A2(net253),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4640_ (.A1(_1407_),
    .A2(net253),
    .B(_2634_),
    .C(net121),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4641_ (.A1(\col_prog_n_reg[275] ),
    .A2(net253),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4642_ (.A1(_1410_),
    .A2(net253),
    .B(_2635_),
    .C(net121),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(\col_prog_n_reg[274] ),
    .A2(net253),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4644_ (.A1(_1413_),
    .A2(net253),
    .B(_2636_),
    .C(net121),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4645_ (.A1(\col_prog_n_reg[273] ),
    .A2(net253),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4646_ (.A1(net324),
    .A2(net253),
    .B(_2637_),
    .C(net121),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4647_ (.A1(\col_prog_n_reg[272] ),
    .A2(net253),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4648_ (.A1(net323),
    .A2(net253),
    .B(_2638_),
    .C(net121),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4649_ (.A1(\col_prog_n_reg[271] ),
    .A2(net253),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4650_ (.A1(_1422_),
    .A2(net253),
    .B(_2639_),
    .C(net121),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4651_ (.A1(\col_prog_n_reg[270] ),
    .A2(net253),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4652_ (.A1(_1425_),
    .A2(net253),
    .B(_2640_),
    .C(net121),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4653_ (.A1(\col_prog_n_reg[269] ),
    .A2(net254),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4654_ (.A1(_1428_),
    .A2(net254),
    .B(_2641_),
    .C(net121),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(\col_prog_n_reg[268] ),
    .A2(net254),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4656_ (.A1(net314),
    .A2(net254),
    .B(_2642_),
    .C(net121),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4657_ (.A1(\col_prog_n_reg[267] ),
    .A2(net254),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4658_ (.A1(net312),
    .A2(net254),
    .B(_2643_),
    .C(net121),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4659_ (.A1(\col_prog_n_reg[266] ),
    .A2(net254),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4660_ (.A1(net310),
    .A2(net254),
    .B(_2644_),
    .C(net121),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4661_ (.A1(\col_prog_n_reg[265] ),
    .A2(net254),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4662_ (.A1(_1440_),
    .A2(net254),
    .B(_2645_),
    .C(net121),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4663_ (.A1(\col_prog_n_reg[264] ),
    .A2(net254),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4664_ (.A1(net306),
    .A2(net254),
    .B(_2646_),
    .C(net121),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4665_ (.A1(\col_prog_n_reg[263] ),
    .A2(_2622_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4666_ (.A1(_1448_),
    .A2(_2622_),
    .B(_2647_),
    .C(_1385_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4667_ (.A1(\col_prog_n_reg[262] ),
    .A2(_2622_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4668_ (.A1(_1451_),
    .A2(_2622_),
    .B(_2648_),
    .C(_1385_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(\col_prog_n_reg[261] ),
    .A2(_2622_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4670_ (.A1(_1454_),
    .A2(_2622_),
    .B(_2649_),
    .C(_1385_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4671_ (.A1(\col_prog_n_reg[260] ),
    .A2(_2622_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4672_ (.A1(_1457_),
    .A2(_2622_),
    .B(_2650_),
    .C(_1385_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4673_ (.A1(\col_prog_n_reg[259] ),
    .A2(_2622_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4674_ (.A1(_1460_),
    .A2(_2622_),
    .B(_2651_),
    .C(_1385_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4675_ (.A1(\col_prog_n_reg[258] ),
    .A2(_2622_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4676_ (.A1(_1463_),
    .A2(_2622_),
    .B(_2652_),
    .C(_1385_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(\col_prog_n_reg[257] ),
    .A2(_2622_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4678_ (.A1(_1466_),
    .A2(_2622_),
    .B(_2653_),
    .C(_1385_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(\col_prog_n_reg[256] ),
    .A2(_2622_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4680_ (.A1(_1469_),
    .A2(_2622_),
    .B(_2654_),
    .C(_1385_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4681_ (.A1(net282),
    .A2(_2297_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(\col_prog_n_reg[255] ),
    .A2(net127),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4683_ (.A1(_1478_),
    .A2(net127),
    .B(_2656_),
    .C(net121),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(\col_prog_n_reg[254] ),
    .A2(net127),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4685_ (.A1(_1481_),
    .A2(net127),
    .B(_2657_),
    .C(net121),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4686_ (.A1(\col_prog_n_reg[253] ),
    .A2(net127),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4687_ (.A1(_1484_),
    .A2(net127),
    .B(_2658_),
    .C(net121),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(\col_prog_n_reg[252] ),
    .A2(net127),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4689_ (.A1(_1487_),
    .A2(net127),
    .B(_2659_),
    .C(net121),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4690_ (.A1(\col_prog_n_reg[251] ),
    .A2(net127),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4691_ (.A1(_1490_),
    .A2(net127),
    .B(_2660_),
    .C(net121),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4692_ (.A1(\col_prog_n_reg[250] ),
    .A2(net127),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4693_ (.A1(_1493_),
    .A2(net127),
    .B(_2661_),
    .C(net121),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4694_ (.A1(\col_prog_n_reg[249] ),
    .A2(net127),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4695_ (.A1(_1392_),
    .A2(net127),
    .B(_2662_),
    .C(net121),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4696_ (.A1(\col_prog_n_reg[248] ),
    .A2(net127),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4697_ (.A1(_1395_),
    .A2(net127),
    .B(_2663_),
    .C(net121),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4698_ (.A1(\col_prog_n_reg[247] ),
    .A2(net127),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4699_ (.A1(_1398_),
    .A2(net127),
    .B(_2664_),
    .C(net121),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4700_ (.A1(\col_prog_n_reg[246] ),
    .A2(net127),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4701_ (.A1(_1401_),
    .A2(net127),
    .B(_2665_),
    .C(net121),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4702_ (.A1(\col_prog_n_reg[245] ),
    .A2(net128),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4703_ (.A1(_1404_),
    .A2(net127),
    .B(_2666_),
    .C(net121),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4704_ (.A1(\col_prog_n_reg[244] ),
    .A2(net128),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4705_ (.A1(_1407_),
    .A2(net128),
    .B(_2667_),
    .C(net121),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4706_ (.A1(\col_prog_n_reg[243] ),
    .A2(net128),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4707_ (.A1(_1410_),
    .A2(net128),
    .B(_2668_),
    .C(net121),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4708_ (.A1(\col_prog_n_reg[242] ),
    .A2(net128),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4709_ (.A1(_1413_),
    .A2(net128),
    .B(_2669_),
    .C(net121),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(\col_prog_n_reg[241] ),
    .A2(net128),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4711_ (.A1(net324),
    .A2(net128),
    .B(_2670_),
    .C(net121),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4712_ (.A1(\col_prog_n_reg[240] ),
    .A2(net128),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4713_ (.A1(net323),
    .A2(net128),
    .B(_2671_),
    .C(net121),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4714_ (.A1(\col_prog_n_reg[239] ),
    .A2(net128),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4715_ (.A1(_1422_),
    .A2(net128),
    .B(_2672_),
    .C(net121),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(\col_prog_n_reg[238] ),
    .A2(net128),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4717_ (.A1(_1425_),
    .A2(net128),
    .B(_2673_),
    .C(net121),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4718_ (.A1(\col_prog_n_reg[237] ),
    .A2(net128),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4719_ (.A1(_1428_),
    .A2(net128),
    .B(_2674_),
    .C(net121),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4720_ (.A1(\col_prog_n_reg[236] ),
    .A2(net128),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4721_ (.A1(net314),
    .A2(_2655_),
    .B(_2675_),
    .C(net121),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(\col_prog_n_reg[235] ),
    .A2(_2655_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4723_ (.A1(net312),
    .A2(_2655_),
    .B(_2676_),
    .C(net121),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4724_ (.A1(\col_prog_n_reg[234] ),
    .A2(_2655_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4725_ (.A1(net310),
    .A2(_2655_),
    .B(_2677_),
    .C(net121),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4726_ (.A1(\col_prog_n_reg[233] ),
    .A2(_2655_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4727_ (.A1(_1440_),
    .A2(_2655_),
    .B(_2678_),
    .C(net121),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(\col_prog_n_reg[232] ),
    .A2(_2655_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4729_ (.A1(net306),
    .A2(_2655_),
    .B(_2679_),
    .C(net121),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4730_ (.A1(net282),
    .A2(\col_prog_n_reg[231] ),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4731_ (.A1(\col_prog_n_reg[231] ),
    .A2(_2298_),
    .B1(_2355_),
    .B2(net268),
    .C(net165),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4732_ (.A1(_2680_),
    .A2(_2681_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4733_ (.A1(net282),
    .A2(\col_prog_n_reg[230] ),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4734_ (.A1(\col_prog_n_reg[230] ),
    .A2(_2298_),
    .B1(_2358_),
    .B2(net268),
    .C(net165),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4735_ (.A1(_2682_),
    .A2(_2683_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4736_ (.A1(net282),
    .A2(\col_prog_n_reg[229] ),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4737_ (.A1(\col_prog_n_reg[229] ),
    .A2(_2298_),
    .B1(_2361_),
    .B2(net268),
    .C(net165),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4738_ (.A1(_2684_),
    .A2(_2685_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4739_ (.A1(net282),
    .A2(\col_prog_n_reg[228] ),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4740_ (.A1(\col_prog_n_reg[228] ),
    .A2(_2298_),
    .B1(_2364_),
    .B2(net268),
    .C(net165),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4741_ (.A1(_2686_),
    .A2(_2687_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4742_ (.A1(net282),
    .A2(\col_prog_n_reg[227] ),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4743_ (.A1(\col_prog_n_reg[227] ),
    .A2(_2298_),
    .B1(_2367_),
    .B2(net268),
    .C(net165),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4744_ (.A1(_2688_),
    .A2(_2689_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4745_ (.A1(net282),
    .A2(\col_prog_n_reg[226] ),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4746_ (.A1(\col_prog_n_reg[226] ),
    .A2(_2298_),
    .B1(_2370_),
    .B2(net268),
    .C(net165),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4747_ (.A1(_2690_),
    .A2(_2691_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4748_ (.A1(net282),
    .A2(\col_prog_n_reg[225] ),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4749_ (.A1(\col_prog_n_reg[225] ),
    .A2(_2298_),
    .B1(_2373_),
    .B2(net268),
    .C(net165),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4750_ (.A1(_2692_),
    .A2(_2693_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4751_ (.A1(net282),
    .A2(\col_prog_n_reg[224] ),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4752_ (.A1(\col_prog_n_reg[224] ),
    .A2(_2298_),
    .B1(_2376_),
    .B2(net268),
    .C(net165),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4753_ (.A1(_2694_),
    .A2(_2695_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4754_ (.A1(\state[3] ),
    .A2(_2300_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4755_ (.A1(\col_prog_n_reg[223] ),
    .A2(net125),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4756_ (.A1(net299),
    .A2(net125),
    .B(_2697_),
    .C(_1385_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(\col_prog_n_reg[222] ),
    .A2(net125),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4758_ (.A1(net297),
    .A2(net125),
    .B(_2698_),
    .C(_1385_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4759_ (.A1(\col_prog_n_reg[221] ),
    .A2(net125),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4760_ (.A1(_1484_),
    .A2(net125),
    .B(_2699_),
    .C(_1385_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4761_ (.A1(\col_prog_n_reg[220] ),
    .A2(net125),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4762_ (.A1(net294),
    .A2(net125),
    .B(_2700_),
    .C(_1385_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(\col_prog_n_reg[219] ),
    .A2(net125),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4764_ (.A1(net291),
    .A2(net125),
    .B(_2701_),
    .C(_1385_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4765_ (.A1(\col_prog_n_reg[218] ),
    .A2(net125),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4766_ (.A1(net289),
    .A2(net125),
    .B(_2702_),
    .C(_1385_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4767_ (.A1(\col_prog_n_reg[217] ),
    .A2(net125),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4768_ (.A1(_1392_),
    .A2(net125),
    .B(_2703_),
    .C(_1385_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4769_ (.A1(\col_prog_n_reg[216] ),
    .A2(net125),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4770_ (.A1(net337),
    .A2(net125),
    .B(_2704_),
    .C(_1385_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(\col_prog_n_reg[215] ),
    .A2(net125),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4772_ (.A1(net335),
    .A2(net125),
    .B(_2705_),
    .C(_1385_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4773_ (.A1(\col_prog_n_reg[214] ),
    .A2(net125),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4774_ (.A1(net333),
    .A2(net125),
    .B(_2706_),
    .C(_1385_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(\col_prog_n_reg[213] ),
    .A2(net126),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4776_ (.A1(_1404_),
    .A2(net126),
    .B(_2707_),
    .C(_1385_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4777_ (.A1(\col_prog_n_reg[212] ),
    .A2(net126),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4778_ (.A1(net330),
    .A2(net126),
    .B(_2708_),
    .C(_1385_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(\col_prog_n_reg[211] ),
    .A2(net126),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4780_ (.A1(net327),
    .A2(net126),
    .B(_2709_),
    .C(_1385_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4781_ (.A1(\col_prog_n_reg[210] ),
    .A2(net126),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4782_ (.A1(net325),
    .A2(net126),
    .B(_2710_),
    .C(_1385_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4783_ (.A1(\col_prog_n_reg[209] ),
    .A2(net126),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4784_ (.A1(net324),
    .A2(net126),
    .B(_2711_),
    .C(_1385_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4785_ (.A1(\col_prog_n_reg[208] ),
    .A2(net126),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4786_ (.A1(net322),
    .A2(net126),
    .B(_2712_),
    .C(_1385_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(\col_prog_n_reg[207] ),
    .A2(net126),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4788_ (.A1(net320),
    .A2(net126),
    .B(_2713_),
    .C(_1385_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4789_ (.A1(\col_prog_n_reg[206] ),
    .A2(_2696_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4790_ (.A1(_1425_),
    .A2(_2696_),
    .B(_2714_),
    .C(_1385_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4791_ (.A1(\col_prog_n_reg[205] ),
    .A2(_2696_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4792_ (.A1(_1428_),
    .A2(_2696_),
    .B(_2715_),
    .C(_1385_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(\col_prog_n_reg[204] ),
    .A2(_2696_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4794_ (.A1(net314),
    .A2(_2696_),
    .B(_2716_),
    .C(_1385_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4795_ (.A1(\col_prog_n_reg[203] ),
    .A2(_2696_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4796_ (.A1(net312),
    .A2(_2696_),
    .B(_2717_),
    .C(_1385_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(\col_prog_n_reg[202] ),
    .A2(_2696_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4798_ (.A1(net310),
    .A2(_2696_),
    .B(_2718_),
    .C(_1385_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4799_ (.A1(\col_prog_n_reg[201] ),
    .A2(_2696_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4800_ (.A1(_1440_),
    .A2(_2696_),
    .B(_2719_),
    .C(_1385_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4801_ (.A1(\col_prog_n_reg[200] ),
    .A2(_2696_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4802_ (.A1(net306),
    .A2(_2696_),
    .B(_2720_),
    .C(_1385_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4803_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[199] ),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4804_ (.A1(\col_prog_n_reg[199] ),
    .A2(_2301_),
    .B1(_2404_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4805_ (.A1(_2721_),
    .A2(_2722_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4806_ (.A1(net282),
    .A2(\col_prog_n_reg[198] ),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4807_ (.A1(\col_prog_n_reg[198] ),
    .A2(_2301_),
    .B1(_2407_),
    .B2(net268),
    .C(net165),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4808_ (.A1(_2723_),
    .A2(_2724_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4809_ (.A1(net282),
    .A2(\col_prog_n_reg[197] ),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4810_ (.A1(\col_prog_n_reg[197] ),
    .A2(_2301_),
    .B1(_2410_),
    .B2(net268),
    .C(net165),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4811_ (.A1(_2725_),
    .A2(_2726_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4812_ (.A1(net282),
    .A2(\col_prog_n_reg[196] ),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4813_ (.A1(\col_prog_n_reg[196] ),
    .A2(_2301_),
    .B1(_2413_),
    .B2(net268),
    .C(net165),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4814_ (.A1(_2727_),
    .A2(_2728_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4815_ (.A1(net282),
    .A2(\col_prog_n_reg[195] ),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4816_ (.A1(\col_prog_n_reg[195] ),
    .A2(_2301_),
    .B1(_2416_),
    .B2(net268),
    .C(net165),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4817_ (.A1(_2729_),
    .A2(_2730_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4818_ (.A1(net282),
    .A2(\col_prog_n_reg[194] ),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4819_ (.A1(\col_prog_n_reg[194] ),
    .A2(_2301_),
    .B1(_2419_),
    .B2(net268),
    .C(net165),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4820_ (.A1(_2731_),
    .A2(_2732_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4821_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[193] ),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4822_ (.A1(\col_prog_n_reg[193] ),
    .A2(_2301_),
    .B1(_2422_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4823_ (.A1(_2733_),
    .A2(_2734_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4824_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[192] ),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4825_ (.A1(\col_prog_n_reg[192] ),
    .A2(_2301_),
    .B1(_2425_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4826_ (.A1(_2735_),
    .A2(_2736_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(\state[3] ),
    .A2(_2303_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4828_ (.A1(\col_prog_n_reg[191] ),
    .A2(net123),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4829_ (.A1(net299),
    .A2(net123),
    .B(_2738_),
    .C(_1385_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4830_ (.A1(\col_prog_n_reg[190] ),
    .A2(net123),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4831_ (.A1(net297),
    .A2(net123),
    .B(_2739_),
    .C(_1385_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(\col_prog_n_reg[189] ),
    .A2(net123),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4833_ (.A1(net295),
    .A2(net123),
    .B(_2740_),
    .C(_1385_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(\col_prog_n_reg[188] ),
    .A2(net123),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4835_ (.A1(net294),
    .A2(net123),
    .B(_2741_),
    .C(_1385_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4836_ (.A1(\col_prog_n_reg[187] ),
    .A2(net123),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4837_ (.A1(net291),
    .A2(net123),
    .B(_2742_),
    .C(_1385_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4838_ (.A1(\col_prog_n_reg[186] ),
    .A2(net123),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4839_ (.A1(net289),
    .A2(net123),
    .B(_2743_),
    .C(_1385_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4840_ (.A1(\col_prog_n_reg[185] ),
    .A2(net123),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4841_ (.A1(net339),
    .A2(net123),
    .B(_2744_),
    .C(_1385_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4842_ (.A1(\col_prog_n_reg[184] ),
    .A2(net123),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4843_ (.A1(net337),
    .A2(net123),
    .B(_2745_),
    .C(_1385_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4844_ (.A1(\col_prog_n_reg[183] ),
    .A2(net123),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4845_ (.A1(net335),
    .A2(net123),
    .B(_2746_),
    .C(_1385_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4846_ (.A1(\col_prog_n_reg[182] ),
    .A2(net123),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4847_ (.A1(net333),
    .A2(net123),
    .B(_2747_),
    .C(_1385_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4848_ (.A1(\col_prog_n_reg[181] ),
    .A2(net124),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4849_ (.A1(net331),
    .A2(net123),
    .B(_2748_),
    .C(_1385_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4850_ (.A1(\col_prog_n_reg[180] ),
    .A2(net124),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4851_ (.A1(net330),
    .A2(net124),
    .B(_2749_),
    .C(_1385_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4852_ (.A1(\col_prog_n_reg[179] ),
    .A2(net124),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4853_ (.A1(net327),
    .A2(net124),
    .B(_2750_),
    .C(_1385_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4854_ (.A1(\col_prog_n_reg[178] ),
    .A2(net124),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4855_ (.A1(net325),
    .A2(net124),
    .B(_2751_),
    .C(_1385_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4856_ (.A1(\col_prog_n_reg[177] ),
    .A2(net124),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4857_ (.A1(net324),
    .A2(net124),
    .B(_2752_),
    .C(_1385_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(\col_prog_n_reg[176] ),
    .A2(net124),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4859_ (.A1(net322),
    .A2(net124),
    .B(_2753_),
    .C(_1385_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4860_ (.A1(\col_prog_n_reg[175] ),
    .A2(net124),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4861_ (.A1(net320),
    .A2(net124),
    .B(_2754_),
    .C(_1385_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4862_ (.A1(\col_prog_n_reg[174] ),
    .A2(_2737_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4863_ (.A1(net318),
    .A2(_2737_),
    .B(_2755_),
    .C(_1385_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(\col_prog_n_reg[173] ),
    .A2(_2737_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4865_ (.A1(net316),
    .A2(_2737_),
    .B(_2756_),
    .C(_1385_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4866_ (.A1(\col_prog_n_reg[172] ),
    .A2(_2737_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4867_ (.A1(net314),
    .A2(_2737_),
    .B(_2757_),
    .C(_1385_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4868_ (.A1(\col_prog_n_reg[171] ),
    .A2(_2737_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4869_ (.A1(net312),
    .A2(_2737_),
    .B(_2758_),
    .C(_1385_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4870_ (.A1(\col_prog_n_reg[170] ),
    .A2(_2737_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4871_ (.A1(net310),
    .A2(_2737_),
    .B(_2759_),
    .C(_1385_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4872_ (.A1(\col_prog_n_reg[169] ),
    .A2(_2737_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4873_ (.A1(_1440_),
    .A2(_2737_),
    .B(_2760_),
    .C(_1385_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(\col_prog_n_reg[168] ),
    .A2(_2737_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4875_ (.A1(net306),
    .A2(_2737_),
    .B(_2761_),
    .C(_1385_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4876_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[167] ),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4877_ (.A1(\col_prog_n_reg[167] ),
    .A2(_2304_),
    .B1(_2453_),
    .B2(net268),
    .C(net166),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4878_ (.A1(_2762_),
    .A2(_2763_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4879_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[166] ),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4880_ (.A1(\col_prog_n_reg[166] ),
    .A2(_2304_),
    .B1(_2456_),
    .B2(net268),
    .C(net166),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4881_ (.A1(_2764_),
    .A2(_2765_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4882_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[165] ),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4883_ (.A1(\col_prog_n_reg[165] ),
    .A2(_2304_),
    .B1(_2459_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4884_ (.A1(_2766_),
    .A2(_2767_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4885_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[164] ),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4886_ (.A1(\col_prog_n_reg[164] ),
    .A2(_2304_),
    .B1(_2462_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4887_ (.A1(_2768_),
    .A2(_2769_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4888_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[163] ),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4889_ (.A1(\col_prog_n_reg[163] ),
    .A2(_2304_),
    .B1(_2465_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4890_ (.A1(_2770_),
    .A2(_2771_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4891_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[162] ),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4892_ (.A1(\col_prog_n_reg[162] ),
    .A2(_2304_),
    .B1(_2468_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4893_ (.A1(_2772_),
    .A2(_2773_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4894_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[161] ),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4895_ (.A1(\col_prog_n_reg[161] ),
    .A2(_2304_),
    .B1(_2471_),
    .B2(net268),
    .C(net166),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4896_ (.A1(_2774_),
    .A2(_2775_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4897_ (.A1(\state[3] ),
    .A2(\col_prog_n_reg[160] ),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4898_ (.A1(\col_prog_n_reg[160] ),
    .A2(_2304_),
    .B1(_2474_),
    .B2(net268),
    .C(_1447_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4899_ (.A1(_2776_),
    .A2(_2777_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4900_ (.A1(\col_prog_n_reg[159] ),
    .A2(_1391_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4901_ (.A1(_1391_),
    .A2(net299),
    .B(_2778_),
    .C(net122),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4902_ (.A1(\col_prog_n_reg[158] ),
    .A2(_1391_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4903_ (.A1(_1391_),
    .A2(net297),
    .B(_2779_),
    .C(net122),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(\col_prog_n_reg[157] ),
    .A2(_1391_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4905_ (.A1(_1391_),
    .A2(net295),
    .B(_2780_),
    .C(net122),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4906_ (.A1(\col_prog_n_reg[156] ),
    .A2(_1391_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4907_ (.A1(_1391_),
    .A2(net294),
    .B(_2781_),
    .C(net122),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4908_ (.A1(\col_prog_n_reg[155] ),
    .A2(_1391_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4909_ (.A1(_1391_),
    .A2(net291),
    .B(_2782_),
    .C(net122),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4910_ (.A1(\col_prog_n_reg[154] ),
    .A2(_1391_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4911_ (.A1(_1391_),
    .A2(net289),
    .B(_2783_),
    .C(net122),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4912_ (.A1(_1447_),
    .A2(_1799_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4913_ (.A1(_1363_),
    .A2(_1683_),
    .B(_1385_),
    .C(_1335_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4914_ (.I(net359),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4915_ (.I(net359),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4916_ (.I(net359),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4917_ (.I(net359),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4918_ (.I(net359),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4919_ (.I(net358),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4920_ (.I(net358),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4921_ (.I(net358),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4922_ (.I(net358),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4923_ (.I(net358),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4924_ (.I(net358),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4925_ (.I(net358),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4926_ (.I(net358),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4927_ (.I(net358),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4928_ (.I(net358),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4929_ (.I(net358),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4930_ (.I(net358),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4931_ (.I(net358),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4932_ (.I(net358),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4933_ (.I(net358),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4934_ (.I(net358),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4935_ (.I(net358),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4936_ (.I(net358),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4937_ (.I(net358),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4938_ (.I(net358),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4939_ (.I(net358),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4940_ (.I(net358),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4941_ (.I(net358),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4942_ (.I(net358),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4943_ (.I(net358),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4944_ (.I(net358),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4945_ (.I(net358),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4946_ (.I(net358),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4947_ (.I(net358),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4948_ (.I(net358),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4949_ (.I(net358),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4950_ (.I(net358),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4951_ (.I(net358),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4952_ (.I(net358),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4953_ (.I(net358),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4954_ (.I(net358),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4955_ (.I(net358),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4956_ (.I(net358),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4957_ (.I(net358),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4958_ (.I(net358),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4959_ (.I(net358),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4960_ (.I(net358),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4961_ (.I(net358),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4962_ (.I(net358),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4963_ (.I(net358),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4964_ (.I(net358),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4965_ (.I(net358),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4966_ (.I(net358),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4967_ (.I(net358),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4968_ (.I(net358),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4969_ (.I(net358),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4970_ (.I(net358),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4971_ (.I(net358),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4972_ (.I(net358),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4973_ (.I(net358),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4974_ (.I(net358),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4975_ (.I(net358),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4976_ (.I(net358),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4977_ (.I(net358),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4978_ (.I(net358),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4979_ (.I(net358),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4980_ (.I(net358),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4981_ (.I(net358),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4982_ (.I(net358),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4983_ (.I(net358),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4984_ (.I(net358),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4985_ (.I(net358),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4986_ (.I(net358),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4987_ (.I(net358),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4988_ (.I(net358),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4989_ (.I(net358),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4990_ (.I(net358),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4991_ (.I(net358),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4992_ (.I(net358),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4993_ (.I(net358),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4994_ (.I(net358),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4995_ (.I(net358),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4996_ (.I(net358),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4997_ (.I(net358),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4998_ (.I(net358),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4999_ (.I(net358),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5000_ (.I(net358),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5001_ (.I(net358),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5002_ (.I(net358),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5003_ (.I(net358),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5004_ (.I(net358),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5005_ (.I(net358),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5006_ (.I(net358),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5007_ (.I(net358),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(net358),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5009_ (.I(net358),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5010_ (.I(net358),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5011_ (.I(net358),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5012_ (.I(net358),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5013_ (.I(net358),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5014_ (.I(net358),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5015_ (.I(net358),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5016_ (.I(net358),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5017_ (.I(net358),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5018_ (.I(net358),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5019_ (.I(net358),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5020_ (.I(net358),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5021_ (.I(net358),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5022_ (.I(net358),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5023_ (.I(net358),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5024_ (.I(net358),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5025_ (.I(net358),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5026_ (.I(net358),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5027_ (.I(net358),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5028_ (.I(net358),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5029_ (.I(net358),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5030_ (.I(net358),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5031_ (.I(net358),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5032_ (.I(net358),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5033_ (.I(net358),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5034_ (.I(net358),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5035_ (.I(net358),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5036_ (.I(net358),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5037_ (.I(net358),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5038_ (.I(net358),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5039_ (.I(net358),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5040_ (.I(net358),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5041_ (.I(net358),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5042_ (.I(net358),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5043_ (.I(net358),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5044_ (.I(net358),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5045_ (.I(net358),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5046_ (.I(net357),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5047_ (.I(net358),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5048_ (.I(net358),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5049_ (.I(net358),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5050_ (.I(net358),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5051_ (.I(net358),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5052_ (.I(net358),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5053_ (.I(net358),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5054_ (.I(net358),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5055_ (.I(net357),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5056_ (.I(net357),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5057_ (.I(net357),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5058_ (.I(net357),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5059_ (.I(net357),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5060_ (.I(net357),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5061_ (.I(net357),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5062_ (.I(net357),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5063_ (.I(net357),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5064_ (.I(net357),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5065_ (.I(net357),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5066_ (.I(net357),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5067_ (.I(net357),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5068_ (.I(net357),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5069_ (.I(net357),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5070_ (.I(net357),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5071_ (.I(net357),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5072_ (.I(net357),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5073_ (.I(net357),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5074_ (.I(net357),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5075_ (.I(net357),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5076_ (.I(net357),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5077_ (.I(net357),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5078_ (.I(net357),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5079_ (.I(net358),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5080_ (.I(net358),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5081_ (.I(net358),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5082_ (.I(net358),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5083_ (.I(net358),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5084_ (.I(net358),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5085_ (.I(net358),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5086_ (.I(net358),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5087_ (.I(net357),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5088_ (.I(net357),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5089_ (.I(net357),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5090_ (.I(net357),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5091_ (.I(net357),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5092_ (.I(net357),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5093_ (.I(net357),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5094_ (.I(net357),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5095_ (.I(net357),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5096_ (.I(net357),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5097_ (.I(net357),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5098_ (.I(net357),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5099_ (.I(net357),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5100_ (.I(net357),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5101_ (.I(net357),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5102_ (.I(net357),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5103_ (.I(net357),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5104_ (.I(net357),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5105_ (.I(net357),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5106_ (.I(net357),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5107_ (.I(net357),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5108_ (.I(net357),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5109_ (.I(net357),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5110_ (.I(net357),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5111_ (.I(net357),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5112_ (.I(net357),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5113_ (.I(net357),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5114_ (.I(net357),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5115_ (.I(net357),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5116_ (.I(net357),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5117_ (.I(net357),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5118_ (.I(net357),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5119_ (.I(net356),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5120_ (.I(net356),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5121_ (.I(net356),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5122_ (.I(net356),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5123_ (.I(net356),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5124_ (.I(net356),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5125_ (.I(net356),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5126_ (.I(net356),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5127_ (.I(net356),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5128_ (.I(net356),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5129_ (.I(net356),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5130_ (.I(net356),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5131_ (.I(net356),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5132_ (.I(net356),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5133_ (.I(net356),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5134_ (.I(net356),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5135_ (.I(net356),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5136_ (.I(net356),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5137_ (.I(net356),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5138_ (.I(net356),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5139_ (.I(net356),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5140_ (.I(net356),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5141_ (.I(net356),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5142_ (.I(net356),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5143_ (.I(net357),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5144_ (.I(net357),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5145_ (.I(net357),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5146_ (.I(net357),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5147_ (.I(net357),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5148_ (.I(net357),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5149_ (.I(net357),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5150_ (.I(net357),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5151_ (.I(net356),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5152_ (.I(net356),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5153_ (.I(net356),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5154_ (.I(net356),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5155_ (.I(net356),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5156_ (.I(net356),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5157_ (.I(net356),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5158_ (.I(net356),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5159_ (.I(net356),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5160_ (.I(net356),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5161_ (.I(net356),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5162_ (.I(net356),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5163_ (.I(net356),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5164_ (.I(net356),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5165_ (.I(net356),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5166_ (.I(net356),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5167_ (.I(net356),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5168_ (.I(net356),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5169_ (.I(net356),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5170_ (.I(net356),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5171_ (.I(net356),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5172_ (.I(net356),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5173_ (.I(net356),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5174_ (.I(net356),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5175_ (.I(net357),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5176_ (.I(net357),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5177_ (.I(net357),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5178_ (.I(net357),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5179_ (.I(net357),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5180_ (.I(net357),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5181_ (.I(net357),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5182_ (.I(net357),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5183_ (.I(net356),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5184_ (.I(net356),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(net356),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5186_ (.I(net356),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5187_ (.I(net356),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5188_ (.I(net356),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5189_ (.I(net356),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5190_ (.I(net356),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5191_ (.I(net356),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5192_ (.I(net356),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5193_ (.I(net356),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5194_ (.I(net356),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5195_ (.I(net356),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5196_ (.I(net356),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5197_ (.I(net356),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5198_ (.I(net356),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5199_ (.I(net356),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5200_ (.I(net356),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5201_ (.I(net356),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5202_ (.I(net356),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5203_ (.I(net356),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5204_ (.I(net356),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5205_ (.I(net356),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5206_ (.I(net356),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5207_ (.I(net357),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5208_ (.I(net357),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5209_ (.I(net357),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5210_ (.I(net357),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5211_ (.I(net357),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5212_ (.I(net357),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5213_ (.I(net357),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5214_ (.I(net357),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5215_ (.I(net356),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5216_ (.I(net356),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5217_ (.I(net356),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5218_ (.I(net356),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5219_ (.I(net356),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5220_ (.I(net356),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5221_ (.I(net356),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5222_ (.I(net356),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5223_ (.I(net356),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5224_ (.I(net356),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5225_ (.I(net356),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5226_ (.I(net356),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5227_ (.I(net356),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5228_ (.I(net356),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5229_ (.I(net356),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5230_ (.I(net356),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5231_ (.I(net356),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5232_ (.I(net356),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5233_ (.I(net356),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5234_ (.I(net356),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5235_ (.I(net356),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5236_ (.I(net356),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5237_ (.I(net356),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5238_ (.I(net356),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5239_ (.I(net357),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5240_ (.I(net357),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5241_ (.I(net357),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5242_ (.I(net357),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5243_ (.I(net357),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5244_ (.I(net357),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5245_ (.I(net357),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5246_ (.I(net357),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5247_ (.I(net356),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5248_ (.I(net356),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5249_ (.I(net356),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5250_ (.I(net356),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5251_ (.I(net356),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5252_ (.I(net356),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5253_ (.I(net356),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5254_ (.I(net356),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5255_ (.I(net356),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5256_ (.I(net356),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5257_ (.I(net356),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5258_ (.I(net356),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5259_ (.I(net356),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5260_ (.I(net356),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5261_ (.I(net356),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5262_ (.I(net356),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5263_ (.I(net356),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5264_ (.I(net356),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5265_ (.I(net356),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5266_ (.I(net356),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5267_ (.I(net356),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5268_ (.I(net356),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5269_ (.I(net356),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5270_ (.I(net356),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5271_ (.I(net359),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5272_ (.I(net359),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5273_ (.I(net359),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5274_ (.I(net359),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5275_ (.I(net359),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5276_ (.I(net358),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5277_ (.I(net358),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5278_ (.I(net358),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5279_ (.I(net358),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5280_ (.I(net358),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5281_ (.I(net358),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5282_ (.I(net357),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5283_ (.I(net356),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5284_ (.I(net357),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5285_ (.I(net356),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5286_ (.I(net356),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5287_ (.I(net359),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5288_ (.I(net359),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5289_ (.I(net359),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5290_ (.I(net358),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5291_ (.I(net359),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5292_ (.I(net359),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5293_ (.I(net359),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5294_ (.I(net359),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5295_ (.I(net359),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5296_ (.I(net358),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5297_ (.I(net358),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5298_ (.I(net358),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5299_ (.I(net358),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5300_ (.I(net358),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5301_ (.I(net357),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5302_ (.I(net357),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5303_ (.I(net356),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5304_ (.I(net356),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5305_ (.I(net356),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5306_ (.I(net356),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5307_ (.I(net357),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5308_ (.I(net357),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5309_ (.I(net357),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5310_ (.I(net357),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5311_ (.I(net357),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5312_ (.I(net357),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5313_ (.I(net356),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5314_ (.I(net356),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5315_ (.I(net356),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5316_ (.I(net357),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5317_ (.I(net356),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5318_ (.I(net357),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5319_ (.I(net356),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5320_ (.I(net356),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5321_ (.I(net356),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5322_ (.I(net356),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5323_ (.I(net356),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5324_ (.I(net357),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5325_ (.I(net356),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5326_ (.I(net356),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5327_ (.I(net356),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5328_ (.I(net357),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5329_ (.I(net357),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5330_ (.I(net357),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5331_ (.I(net356),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5332_ (.I(net357),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5333_ (.I(net357),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5334_ (.I(net356),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5335_ (.I(net357),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5336_ (.I(net356),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5337_ (.I(net356),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5338_ (.I(net356),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5339_ (.I(net359),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5340_ (.I(net358),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5341_ (.I(net358),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5342_ (.I(net358),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5343_ (.I(net358),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5344_ (.I(net358),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5345_ (.I(net358),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5346_ (.I(net358),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5347_ (.I(net358),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5348_ (.I(net358),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5349_ (.I(net358),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5350_ (.I(net44),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5351_ (.I(net359),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5352_ (.I(net44),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5353_ (.I(net44),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5354_ (.I(net359),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5355_ (.I(net359),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5356_ (.I(net359),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5357_ (.I(net359),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5358_ (.I(net359),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5359_ (.I(net359),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5360_ (.I(net359),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5361_ (.I(net44),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5362_ (.I(net359),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5363_ (.I(net359),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5364_ (.I(net359),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5365_ (.I(net359),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5366_ (.I(net44),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5367_ (.I(net359),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5368_ (.I(net44),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5369_ (.I(net44),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5370_ (.I(net359),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5371_ (.I(net359),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5372_ (.I(net359),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5373_ (.I(net359),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5374_ (.I(net359),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5375_ (.I(net359),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5376_ (.I(net359),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5377_ (.I(net44),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5378_ (.I(net359),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5379_ (.I(net359),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5380_ (.I(net359),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(net359),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5382_ (.I(net44),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5383_ (.I(net359),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5384_ (.I(net44),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5385_ (.I(net44),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5386_ (.I(net359),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5387_ (.I(net359),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5388_ (.I(net359),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5389_ (.I(net359),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5390_ (.I(net359),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5391_ (.I(net359),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5392_ (.I(net359),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5393_ (.I(net44),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5394_ (.I(net359),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5395_ (.I(net359),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5396_ (.I(net359),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5397_ (.I(net359),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5398_ (.I(net44),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5399_ (.I(net359),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5400_ (.I(net44),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5401_ (.I(net44),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5402_ (.I(net359),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5403_ (.I(net359),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5404_ (.I(net359),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5405_ (.I(net359),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5406_ (.I(net359),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5407_ (.I(net359),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5408_ (.I(net359),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5409_ (.I(net44),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5410_ (.I(net359),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5411_ (.I(net359),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5412_ (.I(net359),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5413_ (.I(net359),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5414_ (.I(net44),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5415_ (.I(net44),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5416_ (.I(net44),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5417_ (.I(net44),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5418_ (.I(net44),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5419_ (.I(net44),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5420_ (.I(net44),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5421_ (.I(net44),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5422_ (.I(net44),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5423_ (.I(net44),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5424_ (.I(net44),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5425_ (.I(net44),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5426_ (.I(net44),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5427_ (.I(net44),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5428_ (.I(net44),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5429_ (.I(net44),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5430_ (.I(net44),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5431_ (.I(net44),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5432_ (.I(net44),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5433_ (.I(net44),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5434_ (.I(net44),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5435_ (.I(net44),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5436_ (.I(net44),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5437_ (.I(net44),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5438_ (.I(net44),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5439_ (.I(net44),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5440_ (.I(net44),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5441_ (.I(net44),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5442_ (.I(net44),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5443_ (.I(net44),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5444_ (.I(net44),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5445_ (.I(net44),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5446_ (.I(net359),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5447_ (.I(net359),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5448_ (.I(net359),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5449_ (.I(net359),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5450_ (.I(net359),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5451_ (.I(net359),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5452_ (.I(net359),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5453_ (.I(net359),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5454_ (.I(net44),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5455_ (.I(net44),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5456_ (.I(net44),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5457_ (.I(net44),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5458_ (.I(net44),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5459_ (.I(net44),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5460_ (.I(net44),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5461_ (.I(net44),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5462_ (.I(net44),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5463_ (.I(net44),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5464_ (.I(net44),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5465_ (.I(net44),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5466_ (.I(net44),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5467_ (.I(net44),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5468_ (.I(net44),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5469_ (.I(net44),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5470_ (.I(net44),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5471_ (.I(net44),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5472_ (.I(net44),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5473_ (.I(net44),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5474_ (.I(net44),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5475_ (.I(net44),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5476_ (.I(net44),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5477_ (.I(net44),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5478_ (.I(net358),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5479_ (.I(net358),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5480_ (.I(net359),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5481_ (.I(net359),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5482_ (.I(net359),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5483_ (.I(net359),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5484_ (.I(net359),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5485_ (.I(net359),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5486_ (.I(net44),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5487_ (.I(net44),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5488_ (.I(net44),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5489_ (.I(net44),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5490_ (.I(net44),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5491_ (.I(net44),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5492_ (.I(net44),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5493_ (.I(net44),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5494_ (.I(net44),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5495_ (.I(net44),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5496_ (.I(net44),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5497_ (.I(net44),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5498_ (.I(net44),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5499_ (.I(net44),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5500_ (.I(net44),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5501_ (.I(net44),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5502_ (.I(net44),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5503_ (.I(net44),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5504_ (.I(net44),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5505_ (.I(net44),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5506_ (.I(net44),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5507_ (.I(net44),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5508_ (.I(net44),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5509_ (.I(net359),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5510_ (.I(net359),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5511_ (.I(net359),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5512_ (.I(net359),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5513_ (.I(net359),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5514_ (.I(net359),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5515_ (.I(net359),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5516_ (.I(net359),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5517_ (.I(net359),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5518_ (.I(net359),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5519_ (.I(net359),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5520_ (.I(net359),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5521_ (.I(net359),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5522_ (.I(net359),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5523_ (.I(net359),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5524_ (.I(net359),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5525_ (.I(net359),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5526_ (.I(net359),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5527_ (.I(net359),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5528_ (.I(net359),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5529_ (.I(net359),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5530_ (.I(net359),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5531_ (.I(net359),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5532_ (.I(net359),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5533_ (.I(net359),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5534_ (.I(net359),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5535_ (.I(net359),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5536_ (.I(net359),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5537_ (.I(net359),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5538_ (.I(net359),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5539_ (.I(net359),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5540_ (.I(net359),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5541_ (.I(net359),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5542_ (.I(net359),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5543_ (.I(net359),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5544_ (.I(net359),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5545_ (.I(net359),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5546_ (.I(net359),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5547_ (.I(net359),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5548_ (.I(net359),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5549_ (.I(net359),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5550_ (.I(net359),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5551_ (.I(net359),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5552_ (.I(net359),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5553_ (.I(net359),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5554_ (.I(net359),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5555_ (.I(net359),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5556_ (.I(net359),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5557_ (.I(net359),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5558_ (.I(net359),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5559_ (.I(net359),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5560_ (.I(net359),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5561_ (.I(net359),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5562_ (.I(net359),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5563_ (.I(net359),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5564_ (.I(net359),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5565_ (.I(net359),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5566_ (.I(net359),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5567_ (.I(net359),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5568_ (.D(_0658_),
    .SETN(_0003_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\col_prog_n_reg[154] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5569_ (.D(_0659_),
    .SETN(_0004_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\col_prog_n_reg[155] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5570_ (.D(_0660_),
    .SETN(_0005_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[156] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5571_ (.D(_0661_),
    .SETN(_0006_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[157] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5572_ (.D(_0662_),
    .SETN(_0007_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[158] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5573_ (.D(_0663_),
    .SETN(_0008_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[159] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5574_ (.D(_0664_),
    .SETN(_0009_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[160] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5575_ (.D(_0665_),
    .SETN(_0010_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[161] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5576_ (.D(_0666_),
    .SETN(_0011_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[162] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5577_ (.D(_0667_),
    .SETN(_0012_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[163] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5578_ (.D(_0668_),
    .SETN(_0013_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[164] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5579_ (.D(_0669_),
    .SETN(_0014_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[165] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5580_ (.D(_0670_),
    .SETN(_0015_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[166] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5581_ (.D(_0671_),
    .SETN(_0016_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[167] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5582_ (.D(_0672_),
    .SETN(_0017_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[168] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5583_ (.D(_0673_),
    .SETN(_0018_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[169] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5584_ (.D(_0674_),
    .SETN(_0019_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[170] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5585_ (.D(_0675_),
    .SETN(_0020_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\col_prog_n_reg[171] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5586_ (.D(_0676_),
    .SETN(_0021_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\col_prog_n_reg[172] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5587_ (.D(_0677_),
    .SETN(_0022_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\col_prog_n_reg[173] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5588_ (.D(_0678_),
    .SETN(_0023_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\col_prog_n_reg[174] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5589_ (.D(_0679_),
    .SETN(_0024_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[175] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5590_ (.D(_0680_),
    .SETN(_0025_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[176] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5591_ (.D(_0681_),
    .SETN(_0026_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[177] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5592_ (.D(_0682_),
    .SETN(_0027_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\col_prog_n_reg[178] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5593_ (.D(_0683_),
    .SETN(_0028_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\col_prog_n_reg[179] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5594_ (.D(_0684_),
    .SETN(_0029_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[180] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5595_ (.D(_0685_),
    .SETN(_0030_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[181] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5596_ (.D(_0686_),
    .SETN(_0031_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[182] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5597_ (.D(_0687_),
    .SETN(_0032_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[183] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5598_ (.D(_0688_),
    .SETN(_0033_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[184] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5599_ (.D(_0689_),
    .SETN(_0034_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[185] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5600_ (.D(_0690_),
    .SETN(_0035_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[186] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5601_ (.D(_0691_),
    .SETN(_0036_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[187] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5602_ (.D(_0692_),
    .SETN(_0037_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[188] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5603_ (.D(_0693_),
    .SETN(_0038_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[189] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5604_ (.D(_0694_),
    .SETN(_0039_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[190] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5605_ (.D(_0695_),
    .SETN(_0040_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[191] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5606_ (.D(_0696_),
    .SETN(_0041_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[192] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5607_ (.D(_0697_),
    .SETN(_0042_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[193] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5608_ (.D(_0698_),
    .SETN(_0043_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[194] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5609_ (.D(_0699_),
    .SETN(_0044_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[195] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5610_ (.D(_0700_),
    .SETN(_0045_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[196] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5611_ (.D(_0701_),
    .SETN(_0046_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[197] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5612_ (.D(_0702_),
    .SETN(_0047_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[198] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5613_ (.D(_0703_),
    .SETN(_0048_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[199] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5614_ (.D(_0704_),
    .SETN(_0049_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[200] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5615_ (.D(_0705_),
    .SETN(_0050_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[201] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5616_ (.D(_0706_),
    .SETN(_0051_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\col_prog_n_reg[202] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5617_ (.D(_0707_),
    .SETN(_0052_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\col_prog_n_reg[203] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5618_ (.D(_0708_),
    .SETN(_0053_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\col_prog_n_reg[204] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5619_ (.D(_0709_),
    .SETN(_0054_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\col_prog_n_reg[205] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5620_ (.D(_0710_),
    .SETN(_0055_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\col_prog_n_reg[206] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5621_ (.D(_0711_),
    .SETN(_0056_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[207] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5622_ (.D(_0712_),
    .SETN(_0057_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[208] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5623_ (.D(_0713_),
    .SETN(_0058_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\col_prog_n_reg[209] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5624_ (.D(_0714_),
    .SETN(_0059_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\col_prog_n_reg[210] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5625_ (.D(_0715_),
    .SETN(_0060_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\col_prog_n_reg[211] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5626_ (.D(_0716_),
    .SETN(_0061_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[212] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5627_ (.D(_0717_),
    .SETN(_0062_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[213] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5628_ (.D(_0718_),
    .SETN(_0063_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[214] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5629_ (.D(_0719_),
    .SETN(_0064_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\col_prog_n_reg[215] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5630_ (.D(_0720_),
    .SETN(_0065_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[216] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5631_ (.D(_0721_),
    .SETN(_0066_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[217] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5632_ (.D(_0722_),
    .SETN(_0067_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[218] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5633_ (.D(_0723_),
    .SETN(_0068_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\col_prog_n_reg[219] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5634_ (.D(_0724_),
    .SETN(_0069_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[220] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5635_ (.D(_0725_),
    .SETN(_0070_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[221] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5636_ (.D(_0726_),
    .SETN(_0071_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[222] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5637_ (.D(_0727_),
    .SETN(_0072_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\col_prog_n_reg[223] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5638_ (.D(_0728_),
    .SETN(_0073_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[224] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5639_ (.D(_0729_),
    .SETN(_0074_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[225] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5640_ (.D(_0730_),
    .SETN(_0075_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[226] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5641_ (.D(_0731_),
    .SETN(_0076_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[227] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5642_ (.D(_0732_),
    .SETN(_0077_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[228] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5643_ (.D(_0733_),
    .SETN(_0078_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[229] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5644_ (.D(_0734_),
    .SETN(_0079_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[230] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5645_ (.D(_0735_),
    .SETN(_0080_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[231] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5646_ (.D(_0736_),
    .SETN(_0081_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[232] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5647_ (.D(_0737_),
    .SETN(_0082_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[233] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5648_ (.D(_0738_),
    .SETN(_0083_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[234] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5649_ (.D(_0739_),
    .SETN(_0084_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[235] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5650_ (.D(_0740_),
    .SETN(_0085_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\col_prog_n_reg[236] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5651_ (.D(_0741_),
    .SETN(_0086_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\col_prog_n_reg[237] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5652_ (.D(_0742_),
    .SETN(_0087_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\col_prog_n_reg[238] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5653_ (.D(_0743_),
    .SETN(_0088_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\col_prog_n_reg[239] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5654_ (.D(_0744_),
    .SETN(_0089_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\col_prog_n_reg[240] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5655_ (.D(_0745_),
    .SETN(_0090_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[241] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5656_ (.D(_0746_),
    .SETN(_0091_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[242] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5657_ (.D(_0747_),
    .SETN(_0092_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[243] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5658_ (.D(_0748_),
    .SETN(_0093_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[244] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5659_ (.D(_0749_),
    .SETN(_0094_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[245] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5660_ (.D(_0750_),
    .SETN(_0095_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\col_prog_n_reg[246] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5661_ (.D(_0751_),
    .SETN(_0096_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\col_prog_n_reg[247] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5662_ (.D(_0752_),
    .SETN(_0097_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[248] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5663_ (.D(_0753_),
    .SETN(_0098_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[249] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5664_ (.D(_0754_),
    .SETN(_0099_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[250] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5665_ (.D(_0755_),
    .SETN(_0100_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[251] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5666_ (.D(_0756_),
    .SETN(_0101_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[252] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5667_ (.D(_0757_),
    .SETN(_0102_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[253] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5668_ (.D(_0758_),
    .SETN(_0103_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[254] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5669_ (.D(_0759_),
    .SETN(_0104_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[255] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5670_ (.D(_0760_),
    .SETN(_0105_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[256] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5671_ (.D(_0761_),
    .SETN(_0106_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[257] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5672_ (.D(_0762_),
    .SETN(_0107_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[258] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5673_ (.D(_0763_),
    .SETN(_0108_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[259] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5674_ (.D(_0764_),
    .SETN(_0109_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[260] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5675_ (.D(_0765_),
    .SETN(_0110_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\col_prog_n_reg[261] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5676_ (.D(_0766_),
    .SETN(_0111_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[262] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5677_ (.D(_0767_),
    .SETN(_0112_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[263] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5678_ (.D(_0768_),
    .SETN(_0113_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[264] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5679_ (.D(_0769_),
    .SETN(_0114_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[265] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5680_ (.D(_0770_),
    .SETN(_0115_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[266] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5681_ (.D(_0771_),
    .SETN(_0116_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\col_prog_n_reg[267] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5682_ (.D(_0772_),
    .SETN(_0117_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\col_prog_n_reg[268] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5683_ (.D(_0773_),
    .SETN(_0118_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\col_prog_n_reg[269] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5684_ (.D(_0774_),
    .SETN(_0119_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\col_prog_n_reg[270] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5685_ (.D(_0775_),
    .SETN(_0120_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\col_prog_n_reg[271] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5686_ (.D(_0776_),
    .SETN(_0121_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\col_prog_n_reg[272] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5687_ (.D(_0777_),
    .SETN(_0122_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\col_prog_n_reg[273] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5688_ (.D(_0778_),
    .SETN(_0123_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[274] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5689_ (.D(_0779_),
    .SETN(_0124_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[275] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5690_ (.D(_0780_),
    .SETN(_0125_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[276] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5691_ (.D(_0781_),
    .SETN(_0126_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\col_prog_n_reg[277] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5692_ (.D(_0782_),
    .SETN(_0127_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\col_prog_n_reg[278] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5693_ (.D(_0783_),
    .SETN(_0128_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\col_prog_n_reg[279] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5694_ (.D(_0784_),
    .SETN(_0129_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[280] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5695_ (.D(_0785_),
    .SETN(_0130_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[281] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5696_ (.D(_0786_),
    .SETN(_0131_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[282] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5697_ (.D(_0787_),
    .SETN(_0132_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\col_prog_n_reg[283] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5698_ (.D(_0788_),
    .SETN(_0133_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[284] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5699_ (.D(_0789_),
    .SETN(_0134_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[285] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5700_ (.D(_0790_),
    .SETN(_0135_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[286] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5701_ (.D(_0791_),
    .SETN(_0136_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\col_prog_n_reg[287] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5702_ (.D(_0792_),
    .SETN(_0137_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[288] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5703_ (.D(_0793_),
    .SETN(_0138_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[289] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5704_ (.D(_0794_),
    .SETN(_0139_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[290] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5705_ (.D(_0795_),
    .SETN(_0140_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[291] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5706_ (.D(_0796_),
    .SETN(_0141_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[292] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5707_ (.D(_0797_),
    .SETN(_0142_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[293] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5708_ (.D(_0798_),
    .SETN(_0143_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[294] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5709_ (.D(_0799_),
    .SETN(_0144_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[295] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5710_ (.D(_0800_),
    .SETN(_0145_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[296] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5711_ (.D(_0801_),
    .SETN(_0146_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[297] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5712_ (.D(_0802_),
    .SETN(_0147_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[298] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5713_ (.D(_0803_),
    .SETN(_0148_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\col_prog_n_reg[299] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5714_ (.D(_0804_),
    .SETN(_0149_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\col_prog_n_reg[300] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5715_ (.D(_0805_),
    .SETN(_0150_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[301] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5716_ (.D(_0806_),
    .SETN(_0151_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[302] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5717_ (.D(_0807_),
    .SETN(_0152_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[303] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5718_ (.D(_0808_),
    .SETN(_0153_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[304] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5719_ (.D(_0809_),
    .SETN(_0154_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[305] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5720_ (.D(_0810_),
    .SETN(_0155_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[306] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5721_ (.D(_0811_),
    .SETN(_0156_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[307] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5722_ (.D(_0812_),
    .SETN(_0157_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[308] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5723_ (.D(_0813_),
    .SETN(_0158_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\col_prog_n_reg[309] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5724_ (.D(_0814_),
    .SETN(_0159_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[310] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5725_ (.D(_0815_),
    .SETN(_0160_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[311] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5726_ (.D(_0816_),
    .SETN(_0161_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[312] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5727_ (.D(_0817_),
    .SETN(_0162_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[313] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5728_ (.D(_0818_),
    .SETN(_0163_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\col_prog_n_reg[314] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5729_ (.D(_0819_),
    .SETN(_0164_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\col_prog_n_reg[315] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5730_ (.D(_0820_),
    .SETN(_0165_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[316] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5731_ (.D(_0821_),
    .SETN(_0166_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[317] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5732_ (.D(_0822_),
    .SETN(_0167_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[318] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5733_ (.D(_0823_),
    .SETN(_0168_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[319] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5734_ (.D(_0824_),
    .SETN(_0169_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[320] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5735_ (.D(_0825_),
    .SETN(_0170_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[321] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5736_ (.D(_0826_),
    .SETN(_0171_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\col_prog_n_reg[322] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5737_ (.D(_0827_),
    .SETN(_0172_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[323] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5738_ (.D(_0828_),
    .SETN(_0173_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[324] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5739_ (.D(_0829_),
    .SETN(_0174_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\col_prog_n_reg[325] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5740_ (.D(_0830_),
    .SETN(_0175_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[326] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5741_ (.D(_0831_),
    .SETN(_0176_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\col_prog_n_reg[327] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5742_ (.D(_0832_),
    .SETN(_0177_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[328] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5743_ (.D(_0833_),
    .SETN(_0178_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[329] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5744_ (.D(_0834_),
    .SETN(_0179_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[330] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5745_ (.D(_0835_),
    .SETN(_0180_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\col_prog_n_reg[331] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5746_ (.D(_0836_),
    .SETN(_0181_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\col_prog_n_reg[332] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5747_ (.D(_0837_),
    .SETN(_0182_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[333] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5748_ (.D(_0838_),
    .SETN(_0183_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[334] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5749_ (.D(_0839_),
    .SETN(_0184_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\col_prog_n_reg[335] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5750_ (.D(_0840_),
    .SETN(_0185_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\col_prog_n_reg[336] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5751_ (.D(_0841_),
    .SETN(_0186_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[337] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5752_ (.D(_0842_),
    .SETN(_0187_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[338] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5753_ (.D(_0843_),
    .SETN(_0188_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\col_prog_n_reg[339] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5754_ (.D(_0844_),
    .SETN(_0189_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\col_prog_n_reg[340] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5755_ (.D(_0845_),
    .SETN(_0190_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\col_prog_n_reg[341] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5756_ (.D(_0846_),
    .SETN(_0191_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\col_prog_n_reg[342] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5757_ (.D(_0847_),
    .SETN(_0192_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[343] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5758_ (.D(_0848_),
    .SETN(_0193_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[344] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5759_ (.D(_0849_),
    .SETN(_0194_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\col_prog_n_reg[345] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5760_ (.D(_0850_),
    .SETN(_0195_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\col_prog_n_reg[346] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5761_ (.D(_0851_),
    .SETN(_0196_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\col_prog_n_reg[347] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5762_ (.D(_0852_),
    .SETN(_0197_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[348] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5763_ (.D(_0853_),
    .SETN(_0198_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[349] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5764_ (.D(_0854_),
    .SETN(_0199_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\col_prog_n_reg[350] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5765_ (.D(_0855_),
    .SETN(_0200_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\col_prog_n_reg[351] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5766_ (.D(_0856_),
    .SETN(_0201_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[352] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5767_ (.D(_0857_),
    .SETN(_0202_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[353] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5768_ (.D(_0858_),
    .SETN(_0203_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[354] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5769_ (.D(_0859_),
    .SETN(_0204_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[355] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5770_ (.D(_0860_),
    .SETN(_0205_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[356] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5771_ (.D(_0861_),
    .SETN(_0206_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[357] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5772_ (.D(_0862_),
    .SETN(_0207_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[358] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5773_ (.D(_0863_),
    .SETN(_0208_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[359] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5774_ (.D(_0864_),
    .SETN(_0209_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\col_prog_n_reg[360] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5775_ (.D(_0865_),
    .SETN(_0210_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\col_prog_n_reg[361] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5776_ (.D(_0866_),
    .SETN(_0211_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[362] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5777_ (.D(_0867_),
    .SETN(_0212_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[363] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5778_ (.D(_0868_),
    .SETN(_0213_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[364] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5779_ (.D(_0869_),
    .SETN(_0214_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\col_prog_n_reg[365] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5780_ (.D(_0870_),
    .SETN(_0215_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\col_prog_n_reg[366] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5781_ (.D(_0871_),
    .SETN(_0216_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\col_prog_n_reg[367] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5782_ (.D(_0872_),
    .SETN(_0217_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\col_prog_n_reg[368] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5783_ (.D(_0873_),
    .SETN(_0218_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[369] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5784_ (.D(_0874_),
    .SETN(_0219_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\col_prog_n_reg[370] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5785_ (.D(_0875_),
    .SETN(_0220_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[371] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5786_ (.D(_0876_),
    .SETN(_0221_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[372] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5787_ (.D(_0877_),
    .SETN(_0222_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\col_prog_n_reg[373] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5788_ (.D(_0878_),
    .SETN(_0223_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\col_prog_n_reg[374] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5789_ (.D(_0879_),
    .SETN(_0224_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[375] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5790_ (.D(_0880_),
    .SETN(_0225_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[376] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5791_ (.D(_0881_),
    .SETN(_0226_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[377] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5792_ (.D(_0882_),
    .SETN(_0227_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[378] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5793_ (.D(_0883_),
    .SETN(_0228_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\col_prog_n_reg[379] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5794_ (.D(_0884_),
    .SETN(_0229_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\col_prog_n_reg[380] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5795_ (.D(_0885_),
    .SETN(_0230_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\col_prog_n_reg[381] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5796_ (.D(_0886_),
    .SETN(_0231_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\col_prog_n_reg[382] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5797_ (.D(_0887_),
    .SETN(_0232_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\col_prog_n_reg[383] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5798_ (.D(_0888_),
    .SETN(_0233_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[384] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5799_ (.D(_0889_),
    .SETN(_0234_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[385] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5800_ (.D(_0890_),
    .SETN(_0235_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[386] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5801_ (.D(_0891_),
    .SETN(_0236_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[387] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5802_ (.D(_0892_),
    .SETN(_0237_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[388] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5803_ (.D(_0893_),
    .SETN(_0238_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[389] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5804_ (.D(_0894_),
    .SETN(_0239_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[390] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5805_ (.D(_0895_),
    .SETN(_0240_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[391] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5806_ (.D(_0896_),
    .SETN(_0241_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\col_prog_n_reg[392] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5807_ (.D(_0897_),
    .SETN(_0242_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\col_prog_n_reg[393] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5808_ (.D(_0898_),
    .SETN(_0243_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[394] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5809_ (.D(_0899_),
    .SETN(_0244_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[395] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5810_ (.D(_0900_),
    .SETN(_0245_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\col_prog_n_reg[396] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5811_ (.D(_0901_),
    .SETN(_0246_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\col_prog_n_reg[397] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5812_ (.D(_0902_),
    .SETN(_0247_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\col_prog_n_reg[398] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5813_ (.D(_0903_),
    .SETN(_0248_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\col_prog_n_reg[399] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5814_ (.D(_0904_),
    .SETN(_0249_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\col_prog_n_reg[400] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5815_ (.D(_0905_),
    .SETN(_0250_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[401] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5816_ (.D(_0906_),
    .SETN(_0251_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[402] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5817_ (.D(_0907_),
    .SETN(_0252_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[403] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5818_ (.D(_0908_),
    .SETN(_0253_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\col_prog_n_reg[404] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5819_ (.D(_0909_),
    .SETN(_0254_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\col_prog_n_reg[405] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5820_ (.D(_0910_),
    .SETN(_0255_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\col_prog_n_reg[406] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5821_ (.D(_0911_),
    .SETN(_0256_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[407] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5822_ (.D(_0912_),
    .SETN(_0257_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[408] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5823_ (.D(_0913_),
    .SETN(_0258_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[409] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5824_ (.D(_0914_),
    .SETN(_0259_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\col_prog_n_reg[410] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5825_ (.D(_0915_),
    .SETN(_0260_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\col_prog_n_reg[411] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5826_ (.D(_0916_),
    .SETN(_0261_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\col_prog_n_reg[412] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5827_ (.D(_0917_),
    .SETN(_0262_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\col_prog_n_reg[413] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5828_ (.D(_0918_),
    .SETN(_0263_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\col_prog_n_reg[414] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5829_ (.D(_0919_),
    .SETN(_0264_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\col_prog_n_reg[415] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5830_ (.D(_0920_),
    .SETN(_0265_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[416] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5831_ (.D(_0921_),
    .SETN(_0266_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[417] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5832_ (.D(_0922_),
    .SETN(_0267_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[418] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5833_ (.D(_0923_),
    .SETN(_0268_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[419] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5834_ (.D(_0924_),
    .SETN(_0269_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[420] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5835_ (.D(_0925_),
    .SETN(_0270_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[421] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5836_ (.D(_0926_),
    .SETN(_0271_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\col_prog_n_reg[422] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5837_ (.D(_0927_),
    .SETN(_0272_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[423] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5838_ (.D(_0928_),
    .SETN(_0273_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[424] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5839_ (.D(_0929_),
    .SETN(_0274_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[425] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5840_ (.D(_0930_),
    .SETN(_0275_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[426] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5841_ (.D(_0931_),
    .SETN(_0276_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\col_prog_n_reg[427] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5842_ (.D(_0932_),
    .SETN(_0277_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[428] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5843_ (.D(_0933_),
    .SETN(_0278_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[429] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5844_ (.D(_0934_),
    .SETN(_0279_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[430] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5845_ (.D(_0935_),
    .SETN(_0280_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\col_prog_n_reg[431] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5846_ (.D(_0936_),
    .SETN(_0281_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\col_prog_n_reg[432] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5847_ (.D(_0937_),
    .SETN(_0282_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\col_prog_n_reg[433] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5848_ (.D(_0938_),
    .SETN(_0283_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[434] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5849_ (.D(_0939_),
    .SETN(_0284_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[435] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5850_ (.D(_0940_),
    .SETN(_0285_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[436] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5851_ (.D(_0941_),
    .SETN(_0286_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[437] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5852_ (.D(_0942_),
    .SETN(_0287_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[438] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5853_ (.D(_0943_),
    .SETN(_0288_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[439] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5854_ (.D(_0944_),
    .SETN(_0289_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[440] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5855_ (.D(_0945_),
    .SETN(_0290_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[441] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5856_ (.D(_0946_),
    .SETN(_0291_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[442] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5857_ (.D(_0947_),
    .SETN(_0292_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[443] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5858_ (.D(_0948_),
    .SETN(_0293_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[444] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5859_ (.D(_0949_),
    .SETN(_0294_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[445] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5860_ (.D(_0950_),
    .SETN(_0295_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[446] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5861_ (.D(_0951_),
    .SETN(_0296_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[447] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5862_ (.D(_0952_),
    .SETN(_0297_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[448] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5863_ (.D(_0953_),
    .SETN(_0298_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[449] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5864_ (.D(_0954_),
    .SETN(_0299_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[450] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5865_ (.D(_0955_),
    .SETN(_0300_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[451] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5866_ (.D(_0956_),
    .SETN(_0301_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[452] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5867_ (.D(_0957_),
    .SETN(_0302_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[453] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5868_ (.D(_0958_),
    .SETN(_0303_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[454] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5869_ (.D(_0959_),
    .SETN(_0304_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[455] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5870_ (.D(_0960_),
    .SETN(_0305_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[456] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5871_ (.D(_0961_),
    .SETN(_0306_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[457] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5872_ (.D(_0962_),
    .SETN(_0307_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[458] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5873_ (.D(_0963_),
    .SETN(_0308_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[459] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5874_ (.D(_0964_),
    .SETN(_0309_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[460] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5875_ (.D(_0965_),
    .SETN(_0310_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[461] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5876_ (.D(_0966_),
    .SETN(_0311_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[462] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5877_ (.D(_0967_),
    .SETN(_0312_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[463] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5878_ (.D(_0968_),
    .SETN(_0313_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[464] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5879_ (.D(_0969_),
    .SETN(_0314_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\col_prog_n_reg[465] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5880_ (.D(_0970_),
    .SETN(_0315_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[466] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5881_ (.D(_0971_),
    .SETN(_0316_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[467] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5882_ (.D(_0972_),
    .SETN(_0317_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[468] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5883_ (.D(_0973_),
    .SETN(_0318_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[469] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5884_ (.D(_0974_),
    .SETN(_0319_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[470] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5885_ (.D(_0975_),
    .SETN(_0320_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[471] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5886_ (.D(_0976_),
    .SETN(_0321_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[472] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5887_ (.D(_0977_),
    .SETN(_0322_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[473] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5888_ (.D(_0978_),
    .SETN(_0323_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[474] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5889_ (.D(_0979_),
    .SETN(_0324_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[475] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5890_ (.D(_0980_),
    .SETN(_0325_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[476] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5891_ (.D(_0981_),
    .SETN(_0326_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[477] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5892_ (.D(_0982_),
    .SETN(_0327_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[478] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5893_ (.D(_0983_),
    .SETN(_0328_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[479] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5894_ (.D(_0984_),
    .SETN(_0329_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[480] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5895_ (.D(_0985_),
    .SETN(_0330_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[481] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5896_ (.D(_0986_),
    .SETN(_0331_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[482] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5897_ (.D(_0987_),
    .SETN(_0332_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[483] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5898_ (.D(_0988_),
    .SETN(_0333_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\col_prog_n_reg[484] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5899_ (.D(_0989_),
    .SETN(_0334_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\col_prog_n_reg[485] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5900_ (.D(_0990_),
    .SETN(_0335_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[486] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5901_ (.D(_0991_),
    .SETN(_0336_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\col_prog_n_reg[487] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5902_ (.D(_0992_),
    .SETN(_0337_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\col_prog_n_reg[488] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5903_ (.D(_0993_),
    .SETN(_0338_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[489] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5904_ (.D(_0994_),
    .SETN(_0339_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[490] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5905_ (.D(_0995_),
    .SETN(_0340_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\col_prog_n_reg[491] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5906_ (.D(_0996_),
    .SETN(_0341_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\col_prog_n_reg[492] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5907_ (.D(_0997_),
    .SETN(_0342_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[493] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5908_ (.D(_0998_),
    .SETN(_0343_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[494] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5909_ (.D(_0999_),
    .SETN(_0344_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[495] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5910_ (.D(_1000_),
    .SETN(_0345_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\col_prog_n_reg[496] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5911_ (.D(_1001_),
    .SETN(_0346_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\col_prog_n_reg[497] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5912_ (.D(_1002_),
    .SETN(_0347_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[498] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5913_ (.D(_1003_),
    .SETN(_0348_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[499] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5914_ (.D(_1004_),
    .SETN(_0349_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\col_prog_n_reg[500] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5915_ (.D(_1005_),
    .SETN(_0350_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[501] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5916_ (.D(_1006_),
    .SETN(_0351_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[502] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5917_ (.D(_1007_),
    .SETN(_0352_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\col_prog_n_reg[503] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5918_ (.D(_1008_),
    .SETN(_0353_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[504] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5919_ (.D(_1009_),
    .SETN(_0354_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\col_prog_n_reg[505] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5920_ (.D(_1010_),
    .SETN(_0355_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[506] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5921_ (.D(_1011_),
    .SETN(_0356_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\col_prog_n_reg[507] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5922_ (.D(_1012_),
    .SETN(_0357_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[508] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5923_ (.D(_1013_),
    .SETN(_0358_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[509] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5924_ (.D(_1014_),
    .SETN(_0359_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[510] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5925_ (.D(_1015_),
    .SETN(_0360_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\col_prog_n_reg[511] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5926_ (.D(_1016_),
    .SETN(_0361_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\preset_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5927_ (.D(_1017_),
    .SETN(_0362_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\preset_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5928_ (.D(_1018_),
    .SETN(_0363_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\preset_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5929_ (.D(_1019_),
    .SETN(_0364_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\preset_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5930_ (.D(_1020_),
    .SETN(_0365_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\preset_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5931_ (.D(_1021_),
    .SETN(_0366_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\preset_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5932_ (.D(_1022_),
    .SETN(_0367_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\preset_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5933_ (.D(_1023_),
    .SETN(_0368_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\preset_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5934_ (.D(_1024_),
    .SETN(_0369_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\preset_n_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5935_ (.D(_1025_),
    .SETN(_0370_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\preset_n_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5936_ (.D(_1026_),
    .SETN(_0371_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\preset_n_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5937_ (.D(_1027_),
    .SETN(_0372_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\preset_n_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5938_ (.D(_1028_),
    .SETN(_0373_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\preset_n_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5939_ (.D(_1029_),
    .SETN(_0374_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\preset_n_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5940_ (.D(_1030_),
    .SETN(_0375_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\preset_n_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5941_ (.D(_1031_),
    .SETN(_0376_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\preset_n_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _5942_ (.D(_0001_),
    .SETN(_0377_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5943_ (.D(\state[2] ),
    .RN(_0378_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5944_ (.D(_0000_),
    .RN(_0379_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _5945_ (.D(_0002_),
    .RN(_0380_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5946_ (.D(_1032_),
    .RN(_0381_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\sense_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5947_ (.D(_1033_),
    .RN(_0382_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\sense_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5948_ (.D(_1034_),
    .RN(_0383_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\sense_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5949_ (.D(_1035_),
    .RN(_0384_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\sense_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5950_ (.D(_1036_),
    .RN(_0385_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\sense_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5951_ (.D(_1037_),
    .RN(_0386_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\sense_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5952_ (.D(_1038_),
    .RN(_0387_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\sense_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5953_ (.D(_1039_),
    .RN(_0388_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\sense_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5954_ (.D(_1040_),
    .RN(_0389_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\sense_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5955_ (.D(_1041_),
    .RN(_0390_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\sense_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5956_ (.D(_1042_),
    .RN(_0391_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\sense_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5957_ (.D(_1043_),
    .RN(_0392_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\sense_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5958_ (.D(_1044_),
    .RN(_0393_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\sense_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5959_ (.D(_1045_),
    .RN(_0394_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\sense_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5960_ (.D(_1046_),
    .RN(_0395_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\sense_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5961_ (.D(_1047_),
    .RN(_0396_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\sense_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5962_ (.D(_1048_),
    .RN(_0397_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5963_ (.D(_1049_),
    .RN(_0398_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5964_ (.D(_1050_),
    .RN(_0399_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5965_ (.D(_1051_),
    .RN(_0400_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5966_ (.D(_1052_),
    .RN(_0401_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5967_ (.D(_1053_),
    .RN(_0402_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5968_ (.D(_1054_),
    .RN(_0403_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net80));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5969_ (.D(_1055_),
    .RN(_0404_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net81));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5970_ (.D(_1056_),
    .RN(_0405_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net82));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5971_ (.D(_1057_),
    .RN(_0406_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5972_ (.D(_1058_),
    .RN(_0407_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5973_ (.D(_1059_),
    .RN(_0408_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5974_ (.D(_1060_),
    .RN(_0409_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5975_ (.D(_1061_),
    .RN(_0410_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5976_ (.D(_1062_),
    .RN(_0411_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5977_ (.D(_1063_),
    .RN(_0412_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5978_ (.D(_1064_),
    .RN(_0413_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5979_ (.D(_1065_),
    .RN(_0414_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5980_ (.D(_1066_),
    .RN(_0415_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5981_ (.D(_1067_),
    .RN(_0416_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5982_ (.D(_1068_),
    .RN(_0417_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5983_ (.D(_1069_),
    .RN(_0418_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5984_ (.D(_1070_),
    .RN(_0419_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5985_ (.D(_1071_),
    .RN(_0420_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5986_ (.D(_1072_),
    .RN(_0421_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5987_ (.D(_1073_),
    .RN(_0422_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5988_ (.D(_1074_),
    .RN(_0423_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5989_ (.D(_1075_),
    .RN(_0424_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5990_ (.D(_1076_),
    .RN(_0425_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5991_ (.D(_1077_),
    .RN(_0426_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5992_ (.D(_1078_),
    .RN(_0427_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5993_ (.D(_1079_),
    .RN(_0428_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net76));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _5994_ (.D(_1080_),
    .RN(_0429_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5995_ (.D(_1081_),
    .RN(_0430_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5996_ (.D(_1082_),
    .RN(_0431_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5997_ (.D(_1083_),
    .RN(_0432_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5998_ (.D(_1084_),
    .RN(_0433_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5999_ (.D(_1085_),
    .RN(_0434_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6000_ (.D(_1086_),
    .RN(_0435_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6001_ (.D(_1087_),
    .RN(_0436_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6002_ (.D(_1088_),
    .RN(_0437_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6003_ (.D(_1089_),
    .RN(_0438_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6004_ (.D(_1090_),
    .RN(_0439_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6005_ (.D(_1091_),
    .RN(_0440_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6006_ (.D(_1092_),
    .RN(_0441_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6007_ (.D(_1093_),
    .RN(_0442_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6008_ (.D(_1094_),
    .RN(_0443_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\bit_sel_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6009_ (.D(_1095_),
    .RN(_0444_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6010_ (.D(_1096_),
    .RN(_0445_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\bit_sel_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6011_ (.D(_1097_),
    .RN(_0446_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6012_ (.D(_1098_),
    .RN(_0447_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6013_ (.D(_1099_),
    .RN(_0448_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6014_ (.D(_1100_),
    .RN(_0449_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6015_ (.D(_1101_),
    .RN(_0450_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6016_ (.D(_1102_),
    .RN(_0451_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\bit_sel_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6017_ (.D(_1103_),
    .RN(_0452_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\bit_sel_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6018_ (.D(_1104_),
    .RN(_0453_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\bit_sel_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6019_ (.D(_1105_),
    .RN(_0454_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6020_ (.D(_1106_),
    .RN(_0455_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6021_ (.D(_1107_),
    .RN(_0456_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6022_ (.D(_1108_),
    .RN(_0457_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6023_ (.D(_1109_),
    .RN(_0458_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\bit_sel_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6024_ (.D(_1110_),
    .RN(_0459_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6025_ (.D(_1111_),
    .RN(_0460_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\bit_sel_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6026_ (.D(_1112_),
    .RN(_0461_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\bit_sel_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6027_ (.D(_1113_),
    .RN(_0462_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6028_ (.D(_1114_),
    .RN(_0463_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\bit_sel_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6029_ (.D(_1115_),
    .RN(_0464_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6030_ (.D(_1116_),
    .RN(_0465_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6031_ (.D(_1117_),
    .RN(_0466_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6032_ (.D(_1118_),
    .RN(_0467_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\bit_sel_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6033_ (.D(_1119_),
    .RN(_0468_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\bit_sel_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6034_ (.D(_1120_),
    .RN(_0469_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6035_ (.D(_1121_),
    .RN(_0470_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6036_ (.D(_1122_),
    .RN(_0471_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6037_ (.D(_1123_),
    .RN(_0472_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6038_ (.D(_1124_),
    .RN(_0473_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6039_ (.D(_1125_),
    .RN(_0474_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6040_ (.D(_1126_),
    .RN(_0475_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\bit_sel_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6041_ (.D(_1127_),
    .RN(_0476_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6042_ (.D(_1128_),
    .RN(_0477_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6043_ (.D(_1129_),
    .RN(_0478_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6044_ (.D(_1130_),
    .RN(_0479_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6045_ (.D(_1131_),
    .RN(_0480_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6046_ (.D(_1132_),
    .RN(_0481_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\bit_sel_reg[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6047_ (.D(_1133_),
    .RN(_0482_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6048_ (.D(_1134_),
    .RN(_0483_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\bit_sel_reg[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6049_ (.D(_1135_),
    .RN(_0484_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6050_ (.D(_1136_),
    .RN(_0485_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\bit_sel_reg[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6051_ (.D(_1137_),
    .RN(_0486_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\bit_sel_reg[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6052_ (.D(_1138_),
    .RN(_0487_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6053_ (.D(_1139_),
    .RN(_0488_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6054_ (.D(_1140_),
    .RN(_0489_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6055_ (.D(_1141_),
    .RN(_0490_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\bit_sel_reg[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6056_ (.D(_1142_),
    .RN(_0491_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6057_ (.D(_1143_),
    .RN(_0492_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\bit_sel_reg[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6058_ (.D(_1144_),
    .RN(_0493_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6059_ (.D(_1145_),
    .RN(_0494_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\bit_sel_reg[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6060_ (.D(_1146_),
    .RN(_0495_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\bit_sel_reg[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6061_ (.D(_1147_),
    .RN(_0496_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6062_ (.D(_1148_),
    .RN(_0497_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6063_ (.D(_1149_),
    .RN(_0498_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\bit_sel_reg[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6064_ (.D(_1150_),
    .RN(_0499_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\bit_sel_reg[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6065_ (.D(_1151_),
    .RN(_0500_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6066_ (.D(_1152_),
    .RN(_0501_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\bit_sel_reg[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6067_ (.D(_1153_),
    .RN(_0502_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\bit_sel_reg[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6068_ (.D(_1154_),
    .RN(_0503_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\bit_sel_reg[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6069_ (.D(_1155_),
    .SETN(_0504_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\col_prog_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6070_ (.D(_1156_),
    .SETN(_0505_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\col_prog_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6071_ (.D(_1157_),
    .SETN(_0506_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\col_prog_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6072_ (.D(_1158_),
    .SETN(_0507_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\col_prog_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6073_ (.D(_1159_),
    .SETN(_0508_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\col_prog_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6074_ (.D(_1160_),
    .SETN(_0509_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\col_prog_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6075_ (.D(_1161_),
    .SETN(_0510_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\col_prog_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6076_ (.D(_1162_),
    .SETN(_0511_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\col_prog_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6077_ (.D(_1163_),
    .SETN(_0512_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\col_prog_n_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6078_ (.D(_1164_),
    .SETN(_0513_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6079_ (.D(_1165_),
    .SETN(_0514_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6080_ (.D(_1166_),
    .SETN(_0515_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6081_ (.D(_1167_),
    .SETN(_0516_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6082_ (.D(_1168_),
    .SETN(_0517_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6083_ (.D(_1169_),
    .SETN(_0518_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6084_ (.D(_1170_),
    .SETN(_0519_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6085_ (.D(_1171_),
    .SETN(_0520_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6086_ (.D(_1172_),
    .SETN(_0521_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6087_ (.D(_1173_),
    .SETN(_0522_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\col_prog_n_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6088_ (.D(_1174_),
    .SETN(_0523_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6089_ (.D(_1175_),
    .SETN(_0524_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\col_prog_n_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6090_ (.D(_1176_),
    .SETN(_0525_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\col_prog_n_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6091_ (.D(_1177_),
    .SETN(_0526_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6092_ (.D(_1178_),
    .SETN(_0527_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6093_ (.D(_1179_),
    .SETN(_0528_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6094_ (.D(_1180_),
    .SETN(_0529_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6095_ (.D(_1181_),
    .SETN(_0530_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6096_ (.D(_1182_),
    .SETN(_0531_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6097_ (.D(_1183_),
    .SETN(_0532_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6098_ (.D(_1184_),
    .SETN(_0533_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6099_ (.D(_1185_),
    .SETN(_0534_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6100_ (.D(_1186_),
    .SETN(_0535_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6101_ (.D(_1187_),
    .SETN(_0536_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6102_ (.D(_1188_),
    .SETN(_0537_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6103_ (.D(_1189_),
    .SETN(_0538_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6104_ (.D(_1190_),
    .SETN(_0539_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6105_ (.D(_1191_),
    .SETN(_0540_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6106_ (.D(_1192_),
    .SETN(_0541_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6107_ (.D(_1193_),
    .SETN(_0542_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6108_ (.D(_1194_),
    .SETN(_0543_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6109_ (.D(_1195_),
    .SETN(_0544_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6110_ (.D(_1196_),
    .SETN(_0545_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6111_ (.D(_1197_),
    .SETN(_0546_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6112_ (.D(_1198_),
    .SETN(_0547_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6113_ (.D(_1199_),
    .SETN(_0548_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6114_ (.D(_1200_),
    .SETN(_0549_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6115_ (.D(_1201_),
    .SETN(_0550_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6116_ (.D(_1202_),
    .SETN(_0551_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6117_ (.D(_1203_),
    .SETN(_0552_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6118_ (.D(_1204_),
    .SETN(_0553_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6119_ (.D(_1205_),
    .SETN(_0554_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\col_prog_n_reg[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6120_ (.D(_1206_),
    .SETN(_0555_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6121_ (.D(_1207_),
    .SETN(_0556_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\col_prog_n_reg[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6122_ (.D(_1208_),
    .SETN(_0557_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\col_prog_n_reg[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6123_ (.D(_1209_),
    .SETN(_0558_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6124_ (.D(_1210_),
    .SETN(_0559_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6125_ (.D(_1211_),
    .SETN(_0560_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6126_ (.D(_1212_),
    .SETN(_0561_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6127_ (.D(_1213_),
    .SETN(_0562_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6128_ (.D(_1214_),
    .SETN(_0563_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6129_ (.D(_1215_),
    .SETN(_0564_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6130_ (.D(_1216_),
    .SETN(_0565_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6131_ (.D(_1217_),
    .SETN(_0566_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6132_ (.D(_1218_),
    .SETN(_0567_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6133_ (.D(_1219_),
    .SETN(_0568_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6134_ (.D(_1220_),
    .SETN(_0569_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\col_prog_n_reg[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6135_ (.D(_1221_),
    .SETN(_0570_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6136_ (.D(_1222_),
    .SETN(_0571_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6137_ (.D(_1223_),
    .SETN(_0572_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6138_ (.D(_1224_),
    .SETN(_0573_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6139_ (.D(_1225_),
    .SETN(_0574_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6140_ (.D(_1226_),
    .SETN(_0575_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6141_ (.D(_1227_),
    .SETN(_0576_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6142_ (.D(_1228_),
    .SETN(_0577_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6143_ (.D(_1229_),
    .SETN(_0578_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6144_ (.D(_1230_),
    .SETN(_0579_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\col_prog_n_reg[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6145_ (.D(_1231_),
    .SETN(_0580_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6146_ (.D(_1232_),
    .SETN(_0581_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\col_prog_n_reg[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6147_ (.D(_1233_),
    .SETN(_0582_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6148_ (.D(_1234_),
    .SETN(_0583_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6149_ (.D(_1235_),
    .SETN(_0584_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\col_prog_n_reg[80] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6150_ (.D(_1236_),
    .SETN(_0585_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[81] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6151_ (.D(_1237_),
    .SETN(_0586_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[82] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6152_ (.D(_1238_),
    .SETN(_0587_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[83] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6153_ (.D(_1239_),
    .SETN(_0588_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\col_prog_n_reg[84] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6154_ (.D(_1240_),
    .SETN(_0589_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\col_prog_n_reg[85] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6155_ (.D(_1241_),
    .SETN(_0590_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[86] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6156_ (.D(_1242_),
    .SETN(_0591_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\col_prog_n_reg[87] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6157_ (.D(_1243_),
    .SETN(_0592_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[88] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6158_ (.D(_1244_),
    .SETN(_0593_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[89] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6159_ (.D(_1245_),
    .SETN(_0594_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\col_prog_n_reg[90] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6160_ (.D(_1246_),
    .SETN(_0595_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[91] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6161_ (.D(_1247_),
    .SETN(_0596_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\col_prog_n_reg[92] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6162_ (.D(_1248_),
    .SETN(_0597_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[93] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6163_ (.D(_1249_),
    .SETN(_0598_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[94] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6164_ (.D(_1250_),
    .SETN(_0599_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\col_prog_n_reg[95] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6165_ (.D(_1251_),
    .SETN(_0600_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[96] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6166_ (.D(_1252_),
    .SETN(_0601_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[97] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6167_ (.D(_1253_),
    .SETN(_0602_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[98] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6168_ (.D(_1254_),
    .SETN(_0603_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\col_prog_n_reg[99] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6169_ (.D(_1255_),
    .SETN(_0604_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[100] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6170_ (.D(_1256_),
    .SETN(_0605_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[101] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6171_ (.D(_1257_),
    .SETN(_0606_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[102] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6172_ (.D(_1258_),
    .SETN(_0607_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[103] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6173_ (.D(_1259_),
    .SETN(_0608_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[104] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6174_ (.D(_1260_),
    .SETN(_0609_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[105] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6175_ (.D(_1261_),
    .SETN(_0610_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[106] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6176_ (.D(_1262_),
    .SETN(_0611_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\col_prog_n_reg[107] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6177_ (.D(_1263_),
    .SETN(_0612_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\col_prog_n_reg[108] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6178_ (.D(_1264_),
    .SETN(_0613_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\col_prog_n_reg[109] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6179_ (.D(_1265_),
    .SETN(_0614_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\col_prog_n_reg[110] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6180_ (.D(_1266_),
    .SETN(_0615_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\col_prog_n_reg[111] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6181_ (.D(_1267_),
    .SETN(_0616_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\col_prog_n_reg[112] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6182_ (.D(_1268_),
    .SETN(_0617_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\col_prog_n_reg[113] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6183_ (.D(_1269_),
    .SETN(_0618_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\col_prog_n_reg[114] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6184_ (.D(_1270_),
    .SETN(_0619_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[115] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6185_ (.D(_1271_),
    .SETN(_0620_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[116] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6186_ (.D(_1272_),
    .SETN(_0621_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[117] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6187_ (.D(_1273_),
    .SETN(_0622_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[118] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6188_ (.D(_1274_),
    .SETN(_0623_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\col_prog_n_reg[119] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6189_ (.D(_1275_),
    .SETN(_0624_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\col_prog_n_reg[120] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6190_ (.D(_1276_),
    .SETN(_0625_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\col_prog_n_reg[121] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6191_ (.D(_1277_),
    .SETN(_0626_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\col_prog_n_reg[122] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6192_ (.D(_1278_),
    .SETN(_0627_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\col_prog_n_reg[123] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6193_ (.D(_1279_),
    .SETN(_0628_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[124] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6194_ (.D(_1280_),
    .SETN(_0629_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[125] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6195_ (.D(_1281_),
    .SETN(_0630_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[126] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6196_ (.D(_1282_),
    .SETN(_0631_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\col_prog_n_reg[127] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6197_ (.D(_1283_),
    .SETN(_0632_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[128] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6198_ (.D(_1284_),
    .SETN(_0633_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[129] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6199_ (.D(_1285_),
    .SETN(_0634_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[130] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6200_ (.D(_1286_),
    .SETN(_0635_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[131] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6201_ (.D(_1287_),
    .SETN(_0636_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\col_prog_n_reg[132] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6202_ (.D(_1288_),
    .SETN(_0637_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[133] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6203_ (.D(_1289_),
    .SETN(_0638_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\col_prog_n_reg[134] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6204_ (.D(_1290_),
    .SETN(_0639_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\col_prog_n_reg[135] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6205_ (.D(_1291_),
    .SETN(_0640_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[136] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6206_ (.D(_1292_),
    .SETN(_0641_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[137] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6207_ (.D(_1293_),
    .SETN(_0642_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\col_prog_n_reg[138] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6208_ (.D(_1294_),
    .SETN(_0643_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\col_prog_n_reg[139] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6209_ (.D(_1295_),
    .SETN(_0644_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\col_prog_n_reg[140] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6210_ (.D(_1296_),
    .SETN(_0645_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\col_prog_n_reg[141] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6211_ (.D(_1297_),
    .SETN(_0646_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\col_prog_n_reg[142] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6212_ (.D(_1298_),
    .SETN(_0647_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\col_prog_n_reg[143] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6213_ (.D(_1299_),
    .SETN(_0648_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\col_prog_n_reg[144] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6214_ (.D(_1300_),
    .SETN(_0649_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\col_prog_n_reg[145] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6215_ (.D(_1301_),
    .SETN(_0650_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\col_prog_n_reg[146] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6216_ (.D(_1302_),
    .SETN(_0651_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[147] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6217_ (.D(_1303_),
    .SETN(_0652_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[148] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6218_ (.D(_1304_),
    .SETN(_0653_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[149] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6219_ (.D(_1305_),
    .SETN(_0654_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\col_prog_n_reg[150] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6220_ (.D(_1306_),
    .SETN(_0655_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\col_prog_n_reg[151] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6221_ (.D(_1307_),
    .SETN(_0656_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\col_prog_n_reg[152] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6222_ (.D(_1308_),
    .SETN(_0657_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\col_prog_n_reg[153] ));
 efuse_array_64x32 \efuse_gen_depth[0].efuse_array  (.PRESET_N(\preset_n[0] ),
    .SENSE(\sense[0] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[31] ,
    \col_prog_n[30] ,
    \col_prog_n[29] ,
    \col_prog_n[28] ,
    \col_prog_n[27] ,
    \col_prog_n[26] ,
    \col_prog_n[25] ,
    \col_prog_n[24] ,
    \col_prog_n[23] ,
    \col_prog_n[22] ,
    \col_prog_n[21] ,
    \col_prog_n[20] ,
    \col_prog_n[19] ,
    \col_prog_n[18] ,
    \col_prog_n[17] ,
    \col_prog_n[16] ,
    \col_prog_n[15] ,
    \col_prog_n[14] ,
    \col_prog_n[13] ,
    \col_prog_n[12] ,
    \col_prog_n[11] ,
    \col_prog_n[10] ,
    \col_prog_n[9] ,
    \col_prog_n[8] ,
    \col_prog_n[7] ,
    \col_prog_n[6] ,
    \col_prog_n[5] ,
    \col_prog_n[4] ,
    \col_prog_n[3] ,
    \col_prog_n[2] ,
    \col_prog_n[1] ,
    \col_prog_n[0] }),
    .OUT({\efuse_out[31] ,
    \efuse_out[30] ,
    \efuse_out[29] ,
    \efuse_out[28] ,
    \efuse_out[27] ,
    \efuse_out[26] ,
    \efuse_out[25] ,
    \efuse_out[24] ,
    \efuse_out[23] ,
    \efuse_out[22] ,
    \efuse_out[21] ,
    \efuse_out[20] ,
    \efuse_out[19] ,
    \efuse_out[18] ,
    \efuse_out[17] ,
    \efuse_out[16] ,
    \efuse_out[15] ,
    \efuse_out[14] ,
    \efuse_out[13] ,
    \efuse_out[12] ,
    \efuse_out[11] ,
    \efuse_out[10] ,
    \efuse_out[9] ,
    \efuse_out[8] ,
    \efuse_out[7] ,
    \efuse_out[6] ,
    \efuse_out[5] ,
    \efuse_out[4] ,
    \efuse_out[3] ,
    \efuse_out[2] ,
    \efuse_out[1] ,
    \efuse_out[0] }));
 efuse_array_64x32 \efuse_gen_depth[10].efuse_array  (.PRESET_N(\preset_n[10] ),
    .SENSE(\sense[10] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[351] ,
    \col_prog_n[350] ,
    \col_prog_n[349] ,
    \col_prog_n[348] ,
    \col_prog_n[347] ,
    \col_prog_n[346] ,
    \col_prog_n[345] ,
    \col_prog_n[344] ,
    \col_prog_n[343] ,
    \col_prog_n[342] ,
    \col_prog_n[341] ,
    \col_prog_n[340] ,
    \col_prog_n[339] ,
    \col_prog_n[338] ,
    \col_prog_n[337] ,
    \col_prog_n[336] ,
    \col_prog_n[335] ,
    \col_prog_n[334] ,
    \col_prog_n[333] ,
    \col_prog_n[332] ,
    \col_prog_n[331] ,
    \col_prog_n[330] ,
    \col_prog_n[329] ,
    \col_prog_n[328] ,
    \col_prog_n[327] ,
    \col_prog_n[326] ,
    \col_prog_n[325] ,
    \col_prog_n[324] ,
    \col_prog_n[323] ,
    \col_prog_n[322] ,
    \col_prog_n[321] ,
    \col_prog_n[320] }),
    .OUT({\efuse_out[351] ,
    \efuse_out[350] ,
    \efuse_out[349] ,
    \efuse_out[348] ,
    \efuse_out[347] ,
    \efuse_out[346] ,
    \efuse_out[345] ,
    \efuse_out[344] ,
    \efuse_out[343] ,
    \efuse_out[342] ,
    \efuse_out[341] ,
    \efuse_out[340] ,
    \efuse_out[339] ,
    \efuse_out[338] ,
    \efuse_out[337] ,
    \efuse_out[336] ,
    \efuse_out[335] ,
    \efuse_out[334] ,
    \efuse_out[333] ,
    \efuse_out[332] ,
    \efuse_out[331] ,
    \efuse_out[330] ,
    \efuse_out[329] ,
    \efuse_out[328] ,
    \efuse_out[327] ,
    \efuse_out[326] ,
    \efuse_out[325] ,
    \efuse_out[324] ,
    \efuse_out[323] ,
    \efuse_out[322] ,
    \efuse_out[321] ,
    \efuse_out[320] }));
 efuse_array_64x32 \efuse_gen_depth[11].efuse_array  (.PRESET_N(\preset_n[11] ),
    .SENSE(\sense[11] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[383] ,
    \col_prog_n[382] ,
    \col_prog_n[381] ,
    \col_prog_n[380] ,
    \col_prog_n[379] ,
    \col_prog_n[378] ,
    \col_prog_n[377] ,
    \col_prog_n[376] ,
    \col_prog_n[375] ,
    \col_prog_n[374] ,
    \col_prog_n[373] ,
    \col_prog_n[372] ,
    \col_prog_n[371] ,
    \col_prog_n[370] ,
    \col_prog_n[369] ,
    \col_prog_n[368] ,
    \col_prog_n[367] ,
    \col_prog_n[366] ,
    \col_prog_n[365] ,
    \col_prog_n[364] ,
    \col_prog_n[363] ,
    \col_prog_n[362] ,
    \col_prog_n[361] ,
    \col_prog_n[360] ,
    \col_prog_n[359] ,
    \col_prog_n[358] ,
    \col_prog_n[357] ,
    \col_prog_n[356] ,
    \col_prog_n[355] ,
    \col_prog_n[354] ,
    \col_prog_n[353] ,
    \col_prog_n[352] }),
    .OUT({\efuse_out[383] ,
    \efuse_out[382] ,
    \efuse_out[381] ,
    \efuse_out[380] ,
    \efuse_out[379] ,
    \efuse_out[378] ,
    \efuse_out[377] ,
    \efuse_out[376] ,
    \efuse_out[375] ,
    \efuse_out[374] ,
    \efuse_out[373] ,
    \efuse_out[372] ,
    \efuse_out[371] ,
    \efuse_out[370] ,
    \efuse_out[369] ,
    \efuse_out[368] ,
    \efuse_out[367] ,
    \efuse_out[366] ,
    \efuse_out[365] ,
    \efuse_out[364] ,
    \efuse_out[363] ,
    \efuse_out[362] ,
    \efuse_out[361] ,
    \efuse_out[360] ,
    \efuse_out[359] ,
    \efuse_out[358] ,
    \efuse_out[357] ,
    \efuse_out[356] ,
    \efuse_out[355] ,
    \efuse_out[354] ,
    \efuse_out[353] ,
    \efuse_out[352] }));
 efuse_array_64x32 \efuse_gen_depth[12].efuse_array  (.PRESET_N(\preset_n[12] ),
    .SENSE(\sense[12] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[415] ,
    \col_prog_n[414] ,
    \col_prog_n[413] ,
    \col_prog_n[412] ,
    \col_prog_n[411] ,
    \col_prog_n[410] ,
    \col_prog_n[409] ,
    \col_prog_n[408] ,
    \col_prog_n[407] ,
    \col_prog_n[406] ,
    \col_prog_n[405] ,
    \col_prog_n[404] ,
    \col_prog_n[403] ,
    \col_prog_n[402] ,
    \col_prog_n[401] ,
    \col_prog_n[400] ,
    \col_prog_n[399] ,
    \col_prog_n[398] ,
    \col_prog_n[397] ,
    \col_prog_n[396] ,
    \col_prog_n[395] ,
    \col_prog_n[394] ,
    \col_prog_n[393] ,
    \col_prog_n[392] ,
    \col_prog_n[391] ,
    \col_prog_n[390] ,
    \col_prog_n[389] ,
    \col_prog_n[388] ,
    \col_prog_n[387] ,
    \col_prog_n[386] ,
    \col_prog_n[385] ,
    \col_prog_n[384] }),
    .OUT({\efuse_out[415] ,
    \efuse_out[414] ,
    \efuse_out[413] ,
    \efuse_out[412] ,
    \efuse_out[411] ,
    \efuse_out[410] ,
    \efuse_out[409] ,
    \efuse_out[408] ,
    \efuse_out[407] ,
    \efuse_out[406] ,
    \efuse_out[405] ,
    \efuse_out[404] ,
    \efuse_out[403] ,
    \efuse_out[402] ,
    \efuse_out[401] ,
    \efuse_out[400] ,
    \efuse_out[399] ,
    \efuse_out[398] ,
    \efuse_out[397] ,
    \efuse_out[396] ,
    \efuse_out[395] ,
    \efuse_out[394] ,
    \efuse_out[393] ,
    \efuse_out[392] ,
    \efuse_out[391] ,
    \efuse_out[390] ,
    \efuse_out[389] ,
    \efuse_out[388] ,
    \efuse_out[387] ,
    \efuse_out[386] ,
    \efuse_out[385] ,
    \efuse_out[384] }));
 efuse_array_64x32 \efuse_gen_depth[13].efuse_array  (.PRESET_N(\preset_n[13] ),
    .SENSE(\sense[13] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[447] ,
    \col_prog_n[446] ,
    \col_prog_n[445] ,
    \col_prog_n[444] ,
    \col_prog_n[443] ,
    \col_prog_n[442] ,
    \col_prog_n[441] ,
    \col_prog_n[440] ,
    \col_prog_n[439] ,
    \col_prog_n[438] ,
    \col_prog_n[437] ,
    \col_prog_n[436] ,
    \col_prog_n[435] ,
    \col_prog_n[434] ,
    \col_prog_n[433] ,
    \col_prog_n[432] ,
    \col_prog_n[431] ,
    \col_prog_n[430] ,
    \col_prog_n[429] ,
    \col_prog_n[428] ,
    \col_prog_n[427] ,
    \col_prog_n[426] ,
    \col_prog_n[425] ,
    \col_prog_n[424] ,
    \col_prog_n[423] ,
    \col_prog_n[422] ,
    \col_prog_n[421] ,
    \col_prog_n[420] ,
    \col_prog_n[419] ,
    \col_prog_n[418] ,
    \col_prog_n[417] ,
    \col_prog_n[416] }),
    .OUT({\efuse_out[447] ,
    \efuse_out[446] ,
    \efuse_out[445] ,
    \efuse_out[444] ,
    \efuse_out[443] ,
    \efuse_out[442] ,
    \efuse_out[441] ,
    \efuse_out[440] ,
    \efuse_out[439] ,
    \efuse_out[438] ,
    \efuse_out[437] ,
    \efuse_out[436] ,
    \efuse_out[435] ,
    \efuse_out[434] ,
    \efuse_out[433] ,
    \efuse_out[432] ,
    \efuse_out[431] ,
    \efuse_out[430] ,
    \efuse_out[429] ,
    \efuse_out[428] ,
    \efuse_out[427] ,
    \efuse_out[426] ,
    \efuse_out[425] ,
    \efuse_out[424] ,
    \efuse_out[423] ,
    \efuse_out[422] ,
    \efuse_out[421] ,
    \efuse_out[420] ,
    \efuse_out[419] ,
    \efuse_out[418] ,
    \efuse_out[417] ,
    \efuse_out[416] }));
 efuse_array_64x32 \efuse_gen_depth[14].efuse_array  (.PRESET_N(\preset_n[14] ),
    .SENSE(\sense[14] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[479] ,
    \col_prog_n[478] ,
    \col_prog_n[477] ,
    \col_prog_n[476] ,
    \col_prog_n[475] ,
    \col_prog_n[474] ,
    \col_prog_n[473] ,
    \col_prog_n[472] ,
    \col_prog_n[471] ,
    \col_prog_n[470] ,
    \col_prog_n[469] ,
    \col_prog_n[468] ,
    \col_prog_n[467] ,
    \col_prog_n[466] ,
    \col_prog_n[465] ,
    \col_prog_n[464] ,
    \col_prog_n[463] ,
    \col_prog_n[462] ,
    \col_prog_n[461] ,
    \col_prog_n[460] ,
    \col_prog_n[459] ,
    \col_prog_n[458] ,
    \col_prog_n[457] ,
    \col_prog_n[456] ,
    \col_prog_n[455] ,
    \col_prog_n[454] ,
    \col_prog_n[453] ,
    \col_prog_n[452] ,
    \col_prog_n[451] ,
    \col_prog_n[450] ,
    \col_prog_n[449] ,
    \col_prog_n[448] }),
    .OUT({\efuse_out[479] ,
    \efuse_out[478] ,
    \efuse_out[477] ,
    \efuse_out[476] ,
    \efuse_out[475] ,
    \efuse_out[474] ,
    \efuse_out[473] ,
    \efuse_out[472] ,
    \efuse_out[471] ,
    \efuse_out[470] ,
    \efuse_out[469] ,
    \efuse_out[468] ,
    \efuse_out[467] ,
    \efuse_out[466] ,
    \efuse_out[465] ,
    \efuse_out[464] ,
    \efuse_out[463] ,
    \efuse_out[462] ,
    \efuse_out[461] ,
    \efuse_out[460] ,
    \efuse_out[459] ,
    \efuse_out[458] ,
    \efuse_out[457] ,
    \efuse_out[456] ,
    \efuse_out[455] ,
    \efuse_out[454] ,
    \efuse_out[453] ,
    \efuse_out[452] ,
    \efuse_out[451] ,
    \efuse_out[450] ,
    \efuse_out[449] ,
    \efuse_out[448] }));
 efuse_array_64x32 \efuse_gen_depth[15].efuse_array  (.PRESET_N(\preset_n[15] ),
    .SENSE(\sense[15] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[511] ,
    \col_prog_n[510] ,
    \col_prog_n[509] ,
    \col_prog_n[508] ,
    \col_prog_n[507] ,
    \col_prog_n[506] ,
    \col_prog_n[505] ,
    \col_prog_n[504] ,
    \col_prog_n[503] ,
    \col_prog_n[502] ,
    \col_prog_n[501] ,
    \col_prog_n[500] ,
    \col_prog_n[499] ,
    \col_prog_n[498] ,
    \col_prog_n[497] ,
    \col_prog_n[496] ,
    \col_prog_n[495] ,
    \col_prog_n[494] ,
    \col_prog_n[493] ,
    \col_prog_n[492] ,
    \col_prog_n[491] ,
    \col_prog_n[490] ,
    \col_prog_n[489] ,
    \col_prog_n[488] ,
    \col_prog_n[487] ,
    \col_prog_n[486] ,
    \col_prog_n[485] ,
    \col_prog_n[484] ,
    \col_prog_n[483] ,
    \col_prog_n[482] ,
    \col_prog_n[481] ,
    \col_prog_n[480] }),
    .OUT({\efuse_out[511] ,
    \efuse_out[510] ,
    \efuse_out[509] ,
    \efuse_out[508] ,
    \efuse_out[507] ,
    \efuse_out[506] ,
    \efuse_out[505] ,
    \efuse_out[504] ,
    \efuse_out[503] ,
    \efuse_out[502] ,
    \efuse_out[501] ,
    \efuse_out[500] ,
    \efuse_out[499] ,
    \efuse_out[498] ,
    \efuse_out[497] ,
    \efuse_out[496] ,
    \efuse_out[495] ,
    \efuse_out[494] ,
    \efuse_out[493] ,
    \efuse_out[492] ,
    \efuse_out[491] ,
    \efuse_out[490] ,
    \efuse_out[489] ,
    \efuse_out[488] ,
    \efuse_out[487] ,
    \efuse_out[486] ,
    \efuse_out[485] ,
    \efuse_out[484] ,
    \efuse_out[483] ,
    \efuse_out[482] ,
    \efuse_out[481] ,
    \efuse_out[480] }));
 efuse_array_64x32 \efuse_gen_depth[1].efuse_array  (.PRESET_N(\preset_n[1] ),
    .SENSE(\sense[1] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[63] ,
    \col_prog_n[62] ,
    \col_prog_n[61] ,
    \col_prog_n[60] ,
    \col_prog_n[59] ,
    \col_prog_n[58] ,
    \col_prog_n[57] ,
    \col_prog_n[56] ,
    \col_prog_n[55] ,
    \col_prog_n[54] ,
    \col_prog_n[53] ,
    \col_prog_n[52] ,
    \col_prog_n[51] ,
    \col_prog_n[50] ,
    \col_prog_n[49] ,
    \col_prog_n[48] ,
    \col_prog_n[47] ,
    \col_prog_n[46] ,
    \col_prog_n[45] ,
    \col_prog_n[44] ,
    \col_prog_n[43] ,
    \col_prog_n[42] ,
    \col_prog_n[41] ,
    \col_prog_n[40] ,
    \col_prog_n[39] ,
    \col_prog_n[38] ,
    \col_prog_n[37] ,
    \col_prog_n[36] ,
    \col_prog_n[35] ,
    \col_prog_n[34] ,
    \col_prog_n[33] ,
    \col_prog_n[32] }),
    .OUT({\efuse_out[63] ,
    \efuse_out[62] ,
    \efuse_out[61] ,
    \efuse_out[60] ,
    \efuse_out[59] ,
    \efuse_out[58] ,
    \efuse_out[57] ,
    \efuse_out[56] ,
    \efuse_out[55] ,
    \efuse_out[54] ,
    \efuse_out[53] ,
    \efuse_out[52] ,
    \efuse_out[51] ,
    \efuse_out[50] ,
    \efuse_out[49] ,
    \efuse_out[48] ,
    \efuse_out[47] ,
    \efuse_out[46] ,
    \efuse_out[45] ,
    \efuse_out[44] ,
    \efuse_out[43] ,
    \efuse_out[42] ,
    \efuse_out[41] ,
    \efuse_out[40] ,
    \efuse_out[39] ,
    \efuse_out[38] ,
    \efuse_out[37] ,
    \efuse_out[36] ,
    \efuse_out[35] ,
    \efuse_out[34] ,
    \efuse_out[33] ,
    \efuse_out[32] }));
 efuse_array_64x32 \efuse_gen_depth[2].efuse_array  (.PRESET_N(\preset_n[2] ),
    .SENSE(\sense[2] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[95] ,
    \col_prog_n[94] ,
    \col_prog_n[93] ,
    \col_prog_n[92] ,
    \col_prog_n[91] ,
    \col_prog_n[90] ,
    \col_prog_n[89] ,
    \col_prog_n[88] ,
    \col_prog_n[87] ,
    \col_prog_n[86] ,
    \col_prog_n[85] ,
    \col_prog_n[84] ,
    \col_prog_n[83] ,
    \col_prog_n[82] ,
    \col_prog_n[81] ,
    \col_prog_n[80] ,
    \col_prog_n[79] ,
    \col_prog_n[78] ,
    \col_prog_n[77] ,
    \col_prog_n[76] ,
    \col_prog_n[75] ,
    \col_prog_n[74] ,
    \col_prog_n[73] ,
    \col_prog_n[72] ,
    \col_prog_n[71] ,
    \col_prog_n[70] ,
    \col_prog_n[69] ,
    \col_prog_n[68] ,
    \col_prog_n[67] ,
    \col_prog_n[66] ,
    \col_prog_n[65] ,
    \col_prog_n[64] }),
    .OUT({\efuse_out[95] ,
    \efuse_out[94] ,
    \efuse_out[93] ,
    \efuse_out[92] ,
    \efuse_out[91] ,
    \efuse_out[90] ,
    \efuse_out[89] ,
    \efuse_out[88] ,
    \efuse_out[87] ,
    \efuse_out[86] ,
    \efuse_out[85] ,
    \efuse_out[84] ,
    \efuse_out[83] ,
    \efuse_out[82] ,
    \efuse_out[81] ,
    \efuse_out[80] ,
    \efuse_out[79] ,
    \efuse_out[78] ,
    \efuse_out[77] ,
    \efuse_out[76] ,
    \efuse_out[75] ,
    \efuse_out[74] ,
    \efuse_out[73] ,
    \efuse_out[72] ,
    \efuse_out[71] ,
    \efuse_out[70] ,
    \efuse_out[69] ,
    \efuse_out[68] ,
    \efuse_out[67] ,
    \efuse_out[66] ,
    \efuse_out[65] ,
    \efuse_out[64] }));
 efuse_array_64x32 \efuse_gen_depth[3].efuse_array  (.PRESET_N(\preset_n[3] ),
    .SENSE(\sense[3] ),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    net198,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    net206,
    net207,
    \bit_sel[49] ,
    net210,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    net215,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    net224,
    net225,
    \bit_sel[33] ,
    net227,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    net233,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    net242,
    net243,
    \bit_sel[17] ,
    net245,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    net250,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    net219,
    net230,
    \bit_sel[1] ,
    net252}),
    .COL_PROG_N({\col_prog_n[127] ,
    \col_prog_n[126] ,
    \col_prog_n[125] ,
    \col_prog_n[124] ,
    \col_prog_n[123] ,
    \col_prog_n[122] ,
    \col_prog_n[121] ,
    \col_prog_n[120] ,
    \col_prog_n[119] ,
    \col_prog_n[118] ,
    \col_prog_n[117] ,
    \col_prog_n[116] ,
    \col_prog_n[115] ,
    \col_prog_n[114] ,
    \col_prog_n[113] ,
    \col_prog_n[112] ,
    \col_prog_n[111] ,
    \col_prog_n[110] ,
    \col_prog_n[109] ,
    \col_prog_n[108] ,
    \col_prog_n[107] ,
    \col_prog_n[106] ,
    \col_prog_n[105] ,
    \col_prog_n[104] ,
    \col_prog_n[103] ,
    \col_prog_n[102] ,
    \col_prog_n[101] ,
    \col_prog_n[100] ,
    \col_prog_n[99] ,
    \col_prog_n[98] ,
    \col_prog_n[97] ,
    \col_prog_n[96] }),
    .OUT({\efuse_out[127] ,
    \efuse_out[126] ,
    \efuse_out[125] ,
    \efuse_out[124] ,
    \efuse_out[123] ,
    \efuse_out[122] ,
    \efuse_out[121] ,
    \efuse_out[120] ,
    \efuse_out[119] ,
    \efuse_out[118] ,
    \efuse_out[117] ,
    \efuse_out[116] ,
    \efuse_out[115] ,
    \efuse_out[114] ,
    \efuse_out[113] ,
    \efuse_out[112] ,
    \efuse_out[111] ,
    \efuse_out[110] ,
    \efuse_out[109] ,
    \efuse_out[108] ,
    \efuse_out[107] ,
    \efuse_out[106] ,
    \efuse_out[105] ,
    \efuse_out[104] ,
    \efuse_out[103] ,
    \efuse_out[102] ,
    \efuse_out[101] ,
    \efuse_out[100] ,
    \efuse_out[99] ,
    \efuse_out[98] ,
    \efuse_out[97] ,
    \efuse_out[96] }));
 efuse_array_64x32 \efuse_gen_depth[4].efuse_array  (.PRESET_N(\preset_n[4] ),
    .SENSE(\sense[4] ),
    .BIT_SEL({net193,
    net194,
    \bit_sel[61] ,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    \bit_sel[54] ,
    \bit_sel[53] ,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    \bit_sel[38] ,
    \bit_sel[37] ,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    \bit_sel[29] ,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    \bit_sel[22] ,
    \bit_sel[21] ,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    \bit_sel[6] ,
    \bit_sel[5] ,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[159] ,
    \col_prog_n[158] ,
    \col_prog_n[157] ,
    \col_prog_n[156] ,
    \col_prog_n[155] ,
    \col_prog_n[154] ,
    \col_prog_n[153] ,
    \col_prog_n[152] ,
    \col_prog_n[151] ,
    \col_prog_n[150] ,
    \col_prog_n[149] ,
    \col_prog_n[148] ,
    \col_prog_n[147] ,
    \col_prog_n[146] ,
    \col_prog_n[145] ,
    \col_prog_n[144] ,
    \col_prog_n[143] ,
    \col_prog_n[142] ,
    \col_prog_n[141] ,
    \col_prog_n[140] ,
    \col_prog_n[139] ,
    \col_prog_n[138] ,
    \col_prog_n[137] ,
    \col_prog_n[136] ,
    \col_prog_n[135] ,
    \col_prog_n[134] ,
    \col_prog_n[133] ,
    \col_prog_n[132] ,
    \col_prog_n[131] ,
    \col_prog_n[130] ,
    \col_prog_n[129] ,
    \col_prog_n[128] }),
    .OUT({\efuse_out[159] ,
    \efuse_out[158] ,
    \efuse_out[157] ,
    \efuse_out[156] ,
    \efuse_out[155] ,
    \efuse_out[154] ,
    \efuse_out[153] ,
    \efuse_out[152] ,
    \efuse_out[151] ,
    \efuse_out[150] ,
    \efuse_out[149] ,
    \efuse_out[148] ,
    \efuse_out[147] ,
    \efuse_out[146] ,
    \efuse_out[145] ,
    \efuse_out[144] ,
    \efuse_out[143] ,
    \efuse_out[142] ,
    \efuse_out[141] ,
    \efuse_out[140] ,
    \efuse_out[139] ,
    \efuse_out[138] ,
    \efuse_out[137] ,
    \efuse_out[136] ,
    \efuse_out[135] ,
    \efuse_out[134] ,
    \efuse_out[133] ,
    \efuse_out[132] ,
    \efuse_out[131] ,
    \efuse_out[130] ,
    \efuse_out[129] ,
    \efuse_out[128] }));
 efuse_array_64x32 \efuse_gen_depth[5].efuse_array  (.PRESET_N(\preset_n[5] ),
    .SENSE(\sense[5] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[191] ,
    \col_prog_n[190] ,
    \col_prog_n[189] ,
    \col_prog_n[188] ,
    \col_prog_n[187] ,
    \col_prog_n[186] ,
    \col_prog_n[185] ,
    \col_prog_n[184] ,
    \col_prog_n[183] ,
    \col_prog_n[182] ,
    \col_prog_n[181] ,
    \col_prog_n[180] ,
    \col_prog_n[179] ,
    \col_prog_n[178] ,
    \col_prog_n[177] ,
    \col_prog_n[176] ,
    \col_prog_n[175] ,
    \col_prog_n[174] ,
    \col_prog_n[173] ,
    \col_prog_n[172] ,
    \col_prog_n[171] ,
    \col_prog_n[170] ,
    \col_prog_n[169] ,
    \col_prog_n[168] ,
    \col_prog_n[167] ,
    \col_prog_n[166] ,
    \col_prog_n[165] ,
    \col_prog_n[164] ,
    \col_prog_n[163] ,
    \col_prog_n[162] ,
    \col_prog_n[161] ,
    \col_prog_n[160] }),
    .OUT({\efuse_out[191] ,
    \efuse_out[190] ,
    \efuse_out[189] ,
    \efuse_out[188] ,
    \efuse_out[187] ,
    \efuse_out[186] ,
    \efuse_out[185] ,
    \efuse_out[184] ,
    \efuse_out[183] ,
    \efuse_out[182] ,
    \efuse_out[181] ,
    \efuse_out[180] ,
    \efuse_out[179] ,
    \efuse_out[178] ,
    \efuse_out[177] ,
    \efuse_out[176] ,
    \efuse_out[175] ,
    \efuse_out[174] ,
    \efuse_out[173] ,
    \efuse_out[172] ,
    \efuse_out[171] ,
    \efuse_out[170] ,
    \efuse_out[169] ,
    \efuse_out[168] ,
    \efuse_out[167] ,
    \efuse_out[166] ,
    \efuse_out[165] ,
    \efuse_out[164] ,
    \efuse_out[163] ,
    \efuse_out[162] ,
    \efuse_out[161] ,
    \efuse_out[160] }));
 efuse_array_64x32 \efuse_gen_depth[6].efuse_array  (.PRESET_N(\preset_n[6] ),
    .SENSE(\sense[6] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[223] ,
    \col_prog_n[222] ,
    \col_prog_n[221] ,
    \col_prog_n[220] ,
    \col_prog_n[219] ,
    \col_prog_n[218] ,
    \col_prog_n[217] ,
    \col_prog_n[216] ,
    \col_prog_n[215] ,
    \col_prog_n[214] ,
    \col_prog_n[213] ,
    \col_prog_n[212] ,
    \col_prog_n[211] ,
    \col_prog_n[210] ,
    \col_prog_n[209] ,
    \col_prog_n[208] ,
    \col_prog_n[207] ,
    \col_prog_n[206] ,
    \col_prog_n[205] ,
    \col_prog_n[204] ,
    \col_prog_n[203] ,
    \col_prog_n[202] ,
    \col_prog_n[201] ,
    \col_prog_n[200] ,
    \col_prog_n[199] ,
    \col_prog_n[198] ,
    \col_prog_n[197] ,
    \col_prog_n[196] ,
    \col_prog_n[195] ,
    \col_prog_n[194] ,
    \col_prog_n[193] ,
    \col_prog_n[192] }),
    .OUT({\efuse_out[223] ,
    \efuse_out[222] ,
    \efuse_out[221] ,
    \efuse_out[220] ,
    \efuse_out[219] ,
    \efuse_out[218] ,
    \efuse_out[217] ,
    \efuse_out[216] ,
    \efuse_out[215] ,
    \efuse_out[214] ,
    \efuse_out[213] ,
    \efuse_out[212] ,
    \efuse_out[211] ,
    \efuse_out[210] ,
    \efuse_out[209] ,
    \efuse_out[208] ,
    \efuse_out[207] ,
    \efuse_out[206] ,
    \efuse_out[205] ,
    \efuse_out[204] ,
    \efuse_out[203] ,
    \efuse_out[202] ,
    \efuse_out[201] ,
    \efuse_out[200] ,
    \efuse_out[199] ,
    \efuse_out[198] ,
    \efuse_out[197] ,
    \efuse_out[196] ,
    \efuse_out[195] ,
    \efuse_out[194] ,
    \efuse_out[193] ,
    \efuse_out[192] }));
 efuse_array_64x32 \efuse_gen_depth[7].efuse_array  (.PRESET_N(\preset_n[7] ),
    .SENSE(\sense[7] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[255] ,
    \col_prog_n[254] ,
    \col_prog_n[253] ,
    \col_prog_n[252] ,
    \col_prog_n[251] ,
    \col_prog_n[250] ,
    \col_prog_n[249] ,
    \col_prog_n[248] ,
    \col_prog_n[247] ,
    \col_prog_n[246] ,
    \col_prog_n[245] ,
    \col_prog_n[244] ,
    \col_prog_n[243] ,
    \col_prog_n[242] ,
    \col_prog_n[241] ,
    \col_prog_n[240] ,
    \col_prog_n[239] ,
    \col_prog_n[238] ,
    \col_prog_n[237] ,
    \col_prog_n[236] ,
    \col_prog_n[235] ,
    \col_prog_n[234] ,
    \col_prog_n[233] ,
    \col_prog_n[232] ,
    \col_prog_n[231] ,
    \col_prog_n[230] ,
    \col_prog_n[229] ,
    \col_prog_n[228] ,
    \col_prog_n[227] ,
    \col_prog_n[226] ,
    \col_prog_n[225] ,
    \col_prog_n[224] }),
    .OUT({\efuse_out[255] ,
    \efuse_out[254] ,
    \efuse_out[253] ,
    \efuse_out[252] ,
    \efuse_out[251] ,
    \efuse_out[250] ,
    \efuse_out[249] ,
    \efuse_out[248] ,
    \efuse_out[247] ,
    \efuse_out[246] ,
    \efuse_out[245] ,
    \efuse_out[244] ,
    \efuse_out[243] ,
    \efuse_out[242] ,
    \efuse_out[241] ,
    \efuse_out[240] ,
    \efuse_out[239] ,
    \efuse_out[238] ,
    \efuse_out[237] ,
    \efuse_out[236] ,
    \efuse_out[235] ,
    \efuse_out[234] ,
    \efuse_out[233] ,
    \efuse_out[232] ,
    \efuse_out[231] ,
    \efuse_out[230] ,
    \efuse_out[229] ,
    \efuse_out[228] ,
    \efuse_out[227] ,
    \efuse_out[226] ,
    \efuse_out[225] ,
    \efuse_out[224] }));
 efuse_array_64x32 \efuse_gen_depth[8].efuse_array  (.PRESET_N(\preset_n[8] ),
    .SENSE(\sense[8] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[287] ,
    \col_prog_n[286] ,
    \col_prog_n[285] ,
    \col_prog_n[284] ,
    \col_prog_n[283] ,
    \col_prog_n[282] ,
    \col_prog_n[281] ,
    \col_prog_n[280] ,
    \col_prog_n[279] ,
    \col_prog_n[278] ,
    \col_prog_n[277] ,
    \col_prog_n[276] ,
    \col_prog_n[275] ,
    \col_prog_n[274] ,
    \col_prog_n[273] ,
    \col_prog_n[272] ,
    \col_prog_n[271] ,
    \col_prog_n[270] ,
    \col_prog_n[269] ,
    \col_prog_n[268] ,
    \col_prog_n[267] ,
    \col_prog_n[266] ,
    \col_prog_n[265] ,
    \col_prog_n[264] ,
    \col_prog_n[263] ,
    \col_prog_n[262] ,
    \col_prog_n[261] ,
    \col_prog_n[260] ,
    \col_prog_n[259] ,
    \col_prog_n[258] ,
    \col_prog_n[257] ,
    \col_prog_n[256] }),
    .OUT({\efuse_out[287] ,
    \efuse_out[286] ,
    \efuse_out[285] ,
    \efuse_out[284] ,
    \efuse_out[283] ,
    \efuse_out[282] ,
    \efuse_out[281] ,
    \efuse_out[280] ,
    \efuse_out[279] ,
    \efuse_out[278] ,
    \efuse_out[277] ,
    \efuse_out[276] ,
    \efuse_out[275] ,
    \efuse_out[274] ,
    \efuse_out[273] ,
    \efuse_out[272] ,
    \efuse_out[271] ,
    \efuse_out[270] ,
    \efuse_out[269] ,
    \efuse_out[268] ,
    \efuse_out[267] ,
    \efuse_out[266] ,
    \efuse_out[265] ,
    \efuse_out[264] ,
    \efuse_out[263] ,
    \efuse_out[262] ,
    \efuse_out[261] ,
    \efuse_out[260] ,
    \efuse_out[259] ,
    \efuse_out[258] ,
    \efuse_out[257] ,
    \efuse_out[256] }));
 efuse_array_64x32 \efuse_gen_depth[9].efuse_array  (.PRESET_N(\preset_n[9] ),
    .SENSE(\sense[9] ),
    .BIT_SEL({net193,
    net194,
    net195,
    net196,
    net198,
    net199,
    net200,
    net201,
    net202,
    net203,
    net204,
    net205,
    net206,
    net207,
    net209,
    net210,
    net211,
    net212,
    net213,
    net214,
    net215,
    net216,
    net217,
    net218,
    net220,
    net221,
    net222,
    net223,
    net224,
    net225,
    net226,
    net227,
    net228,
    net229,
    net231,
    net232,
    net233,
    net234,
    net235,
    net236,
    net237,
    net238,
    net239,
    net240,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net189,
    net190,
    net191,
    net192,
    net197,
    net208,
    net219,
    net230,
    net241,
    net252}),
    .COL_PROG_N({\col_prog_n[319] ,
    \col_prog_n[318] ,
    \col_prog_n[317] ,
    \col_prog_n[316] ,
    \col_prog_n[315] ,
    \col_prog_n[314] ,
    \col_prog_n[313] ,
    \col_prog_n[312] ,
    \col_prog_n[311] ,
    \col_prog_n[310] ,
    \col_prog_n[309] ,
    \col_prog_n[308] ,
    \col_prog_n[307] ,
    \col_prog_n[306] ,
    \col_prog_n[305] ,
    \col_prog_n[304] ,
    \col_prog_n[303] ,
    \col_prog_n[302] ,
    \col_prog_n[301] ,
    \col_prog_n[300] ,
    \col_prog_n[299] ,
    \col_prog_n[298] ,
    \col_prog_n[297] ,
    \col_prog_n[296] ,
    \col_prog_n[295] ,
    \col_prog_n[294] ,
    \col_prog_n[293] ,
    \col_prog_n[292] ,
    \col_prog_n[291] ,
    \col_prog_n[290] ,
    \col_prog_n[289] ,
    \col_prog_n[288] }),
    .OUT({\efuse_out[319] ,
    \efuse_out[318] ,
    \efuse_out[317] ,
    \efuse_out[316] ,
    \efuse_out[315] ,
    \efuse_out[314] ,
    \efuse_out[313] ,
    \efuse_out[312] ,
    \efuse_out[311] ,
    \efuse_out[310] ,
    \efuse_out[309] ,
    \efuse_out[308] ,
    \efuse_out[307] ,
    \efuse_out[306] ,
    \efuse_out[305] ,
    \efuse_out[304] ,
    \efuse_out[303] ,
    \efuse_out[302] ,
    \efuse_out[301] ,
    \efuse_out[300] ,
    \efuse_out[299] ,
    \efuse_out[298] ,
    \efuse_out[297] ,
    \efuse_out[296] ,
    \efuse_out[295] ,
    \efuse_out[294] ,
    \efuse_out[293] ,
    \efuse_out[292] ,
    \efuse_out[291] ,
    \efuse_out[290] ,
    \efuse_out[289] ,
    \efuse_out[288] }));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[0].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[0] ),
    .S(write_enable_i),
    .Z(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[100].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[100] ),
    .S(write_enable_i),
    .Z(\col_prog_n[100] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[101].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[101] ),
    .S(write_enable_i),
    .Z(\col_prog_n[101] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[102].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[102] ),
    .S(write_enable_i),
    .Z(\col_prog_n[102] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[103].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[103] ),
    .S(write_enable_i),
    .Z(\col_prog_n[103] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[104].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[104] ),
    .S(write_enable_i),
    .Z(\col_prog_n[104] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[105].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[105] ),
    .S(write_enable_i),
    .Z(\col_prog_n[105] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[106].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[106] ),
    .S(write_enable_i),
    .Z(\col_prog_n[106] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[107].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[107] ),
    .S(write_enable_i),
    .Z(\col_prog_n[107] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[108].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[108] ),
    .S(write_enable_i),
    .Z(\col_prog_n[108] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[109].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[109] ),
    .S(write_enable_i),
    .Z(\col_prog_n[109] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[10].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[10] ),
    .S(write_enable_i),
    .Z(\col_prog_n[10] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[110].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[110] ),
    .S(write_enable_i),
    .Z(\col_prog_n[110] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[111].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[111] ),
    .S(write_enable_i),
    .Z(\col_prog_n[111] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[112].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[112] ),
    .S(write_enable_i),
    .Z(\col_prog_n[112] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[113].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[113] ),
    .S(write_enable_i),
    .Z(\col_prog_n[113] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[114].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[114] ),
    .S(write_enable_i),
    .Z(\col_prog_n[114] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[115].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[115] ),
    .S(write_enable_i),
    .Z(\col_prog_n[115] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[116].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[116] ),
    .S(write_enable_i),
    .Z(\col_prog_n[116] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[117].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[117] ),
    .S(write_enable_i),
    .Z(\col_prog_n[117] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[118].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[118] ),
    .S(write_enable_i),
    .Z(\col_prog_n[118] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[119].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[119] ),
    .S(write_enable_i),
    .Z(\col_prog_n[119] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[11].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[11] ),
    .S(write_enable_i),
    .Z(\col_prog_n[11] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[120].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[120] ),
    .S(write_enable_i),
    .Z(\col_prog_n[120] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[121].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[121] ),
    .S(write_enable_i),
    .Z(\col_prog_n[121] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[122].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[122] ),
    .S(write_enable_i),
    .Z(\col_prog_n[122] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[123].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[123] ),
    .S(write_enable_i),
    .Z(\col_prog_n[123] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[124].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[124] ),
    .S(write_enable_i),
    .Z(\col_prog_n[124] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[125].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[125] ),
    .S(write_enable_i),
    .Z(\col_prog_n[125] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[126].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[126] ),
    .S(write_enable_i),
    .Z(\col_prog_n[126] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[127].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[127] ),
    .S(write_enable_i),
    .Z(\col_prog_n[127] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[128].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[128] ),
    .S(write_enable_i),
    .Z(\col_prog_n[128] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[129].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[129] ),
    .S(write_enable_i),
    .Z(\col_prog_n[129] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[12].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[12] ),
    .S(write_enable_i),
    .Z(\col_prog_n[12] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[130].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[130] ),
    .S(write_enable_i),
    .Z(\col_prog_n[130] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[131].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[131] ),
    .S(write_enable_i),
    .Z(\col_prog_n[131] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[132].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[132] ),
    .S(write_enable_i),
    .Z(\col_prog_n[132] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[133].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[133] ),
    .S(write_enable_i),
    .Z(\col_prog_n[133] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[134].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[134] ),
    .S(write_enable_i),
    .Z(\col_prog_n[134] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[135].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[135] ),
    .S(write_enable_i),
    .Z(\col_prog_n[135] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[136].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[136] ),
    .S(write_enable_i),
    .Z(\col_prog_n[136] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[137].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[137] ),
    .S(write_enable_i),
    .Z(\col_prog_n[137] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[138].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[138] ),
    .S(write_enable_i),
    .Z(\col_prog_n[138] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[139].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[139] ),
    .S(write_enable_i),
    .Z(\col_prog_n[139] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[13].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[13] ),
    .S(write_enable_i),
    .Z(\col_prog_n[13] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[140].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[140] ),
    .S(write_enable_i),
    .Z(\col_prog_n[140] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[141].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[141] ),
    .S(write_enable_i),
    .Z(\col_prog_n[141] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[142].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[142] ),
    .S(write_enable_i),
    .Z(\col_prog_n[142] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[143].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[143] ),
    .S(write_enable_i),
    .Z(\col_prog_n[143] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[144].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[144] ),
    .S(write_enable_i),
    .Z(\col_prog_n[144] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[145].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[145] ),
    .S(write_enable_i),
    .Z(\col_prog_n[145] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[146].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[146] ),
    .S(write_enable_i),
    .Z(\col_prog_n[146] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[147].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[147] ),
    .S(write_enable_i),
    .Z(\col_prog_n[147] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[148].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[148] ),
    .S(write_enable_i),
    .Z(\col_prog_n[148] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[149].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[149] ),
    .S(write_enable_i),
    .Z(\col_prog_n[149] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[14].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[14] ),
    .S(write_enable_i),
    .Z(\col_prog_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[150].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[150] ),
    .S(write_enable_i),
    .Z(\col_prog_n[150] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[151].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[151] ),
    .S(write_enable_i),
    .Z(\col_prog_n[151] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[152].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[152] ),
    .S(write_enable_i),
    .Z(\col_prog_n[152] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[153].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[153] ),
    .S(write_enable_i),
    .Z(\col_prog_n[153] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[154].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[154] ),
    .S(write_enable_i),
    .Z(\col_prog_n[154] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[155].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[155] ),
    .S(write_enable_i),
    .Z(\col_prog_n[155] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[156].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[156] ),
    .S(write_enable_i),
    .Z(\col_prog_n[156] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[157].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[157] ),
    .S(write_enable_i),
    .Z(\col_prog_n[157] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[158].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[158] ),
    .S(write_enable_i),
    .Z(\col_prog_n[158] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[159].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[159] ),
    .S(write_enable_i),
    .Z(\col_prog_n[159] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[15].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[15] ),
    .S(write_enable_i),
    .Z(\col_prog_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[160].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[160] ),
    .S(write_enable_i),
    .Z(\col_prog_n[160] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[161].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[161] ),
    .S(write_enable_i),
    .Z(\col_prog_n[161] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[162].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[162] ),
    .S(write_enable_i),
    .Z(\col_prog_n[162] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[163].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[163] ),
    .S(write_enable_i),
    .Z(\col_prog_n[163] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[164].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[164] ),
    .S(write_enable_i),
    .Z(\col_prog_n[164] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[165].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[165] ),
    .S(write_enable_i),
    .Z(\col_prog_n[165] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[166].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[166] ),
    .S(write_enable_i),
    .Z(\col_prog_n[166] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[167].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[167] ),
    .S(write_enable_i),
    .Z(\col_prog_n[167] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[168].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[168] ),
    .S(write_enable_i),
    .Z(\col_prog_n[168] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[169].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[169] ),
    .S(write_enable_i),
    .Z(\col_prog_n[169] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[16].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[16] ),
    .S(write_enable_i),
    .Z(\col_prog_n[16] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[170].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[170] ),
    .S(write_enable_i),
    .Z(\col_prog_n[170] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[171].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[171] ),
    .S(write_enable_i),
    .Z(\col_prog_n[171] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[172].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[172] ),
    .S(write_enable_i),
    .Z(\col_prog_n[172] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[173].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[173] ),
    .S(write_enable_i),
    .Z(\col_prog_n[173] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[174].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[174] ),
    .S(write_enable_i),
    .Z(\col_prog_n[174] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[175].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[175] ),
    .S(write_enable_i),
    .Z(\col_prog_n[175] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[176].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[176] ),
    .S(write_enable_i),
    .Z(\col_prog_n[176] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[177].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[177] ),
    .S(write_enable_i),
    .Z(\col_prog_n[177] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[178].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[178] ),
    .S(write_enable_i),
    .Z(\col_prog_n[178] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[179].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[179] ),
    .S(write_enable_i),
    .Z(\col_prog_n[179] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[17].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[17] ),
    .S(write_enable_i),
    .Z(\col_prog_n[17] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[180].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[180] ),
    .S(write_enable_i),
    .Z(\col_prog_n[180] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[181].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[181] ),
    .S(write_enable_i),
    .Z(\col_prog_n[181] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[182].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[182] ),
    .S(write_enable_i),
    .Z(\col_prog_n[182] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[183].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[183] ),
    .S(write_enable_i),
    .Z(\col_prog_n[183] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[184].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[184] ),
    .S(write_enable_i),
    .Z(\col_prog_n[184] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[185].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[185] ),
    .S(write_enable_i),
    .Z(\col_prog_n[185] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[186].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[186] ),
    .S(write_enable_i),
    .Z(\col_prog_n[186] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[187].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[187] ),
    .S(write_enable_i),
    .Z(\col_prog_n[187] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[188].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[188] ),
    .S(write_enable_i),
    .Z(\col_prog_n[188] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[189].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[189] ),
    .S(write_enable_i),
    .Z(\col_prog_n[189] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[18].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[18] ),
    .S(write_enable_i),
    .Z(\col_prog_n[18] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[190].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[190] ),
    .S(write_enable_i),
    .Z(\col_prog_n[190] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[191].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[191] ),
    .S(write_enable_i),
    .Z(\col_prog_n[191] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[192].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[192] ),
    .S(write_enable_i),
    .Z(\col_prog_n[192] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[193].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[193] ),
    .S(write_enable_i),
    .Z(\col_prog_n[193] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[194].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[194] ),
    .S(write_enable_i),
    .Z(\col_prog_n[194] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[195].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[195] ),
    .S(write_enable_i),
    .Z(\col_prog_n[195] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[196].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[196] ),
    .S(write_enable_i),
    .Z(\col_prog_n[196] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[197].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[197] ),
    .S(write_enable_i),
    .Z(\col_prog_n[197] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[198].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[198] ),
    .S(write_enable_i),
    .Z(\col_prog_n[198] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[199].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[199] ),
    .S(write_enable_i),
    .Z(\col_prog_n[199] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[19].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[19] ),
    .S(write_enable_i),
    .Z(\col_prog_n[19] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[1].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[1] ),
    .S(write_enable_i),
    .Z(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[200].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[200] ),
    .S(write_enable_i),
    .Z(\col_prog_n[200] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[201].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[201] ),
    .S(write_enable_i),
    .Z(\col_prog_n[201] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[202].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[202] ),
    .S(write_enable_i),
    .Z(\col_prog_n[202] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[203].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[203] ),
    .S(write_enable_i),
    .Z(\col_prog_n[203] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[204].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[204] ),
    .S(write_enable_i),
    .Z(\col_prog_n[204] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[205].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[205] ),
    .S(write_enable_i),
    .Z(\col_prog_n[205] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[206].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[206] ),
    .S(write_enable_i),
    .Z(\col_prog_n[206] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[207].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[207] ),
    .S(write_enable_i),
    .Z(\col_prog_n[207] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[208].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[208] ),
    .S(write_enable_i),
    .Z(\col_prog_n[208] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[209].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[209] ),
    .S(write_enable_i),
    .Z(\col_prog_n[209] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[20].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[20] ),
    .S(write_enable_i),
    .Z(\col_prog_n[20] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[210].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[210] ),
    .S(write_enable_i),
    .Z(\col_prog_n[210] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[211].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[211] ),
    .S(write_enable_i),
    .Z(\col_prog_n[211] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[212].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[212] ),
    .S(write_enable_i),
    .Z(\col_prog_n[212] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[213].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[213] ),
    .S(write_enable_i),
    .Z(\col_prog_n[213] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[214].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[214] ),
    .S(write_enable_i),
    .Z(\col_prog_n[214] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[215].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[215] ),
    .S(write_enable_i),
    .Z(\col_prog_n[215] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[216].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[216] ),
    .S(write_enable_i),
    .Z(\col_prog_n[216] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[217].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[217] ),
    .S(write_enable_i),
    .Z(\col_prog_n[217] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[218].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[218] ),
    .S(write_enable_i),
    .Z(\col_prog_n[218] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[219].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[219] ),
    .S(write_enable_i),
    .Z(\col_prog_n[219] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[21].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[21] ),
    .S(write_enable_i),
    .Z(\col_prog_n[21] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[220].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[220] ),
    .S(write_enable_i),
    .Z(\col_prog_n[220] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[221].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[221] ),
    .S(write_enable_i),
    .Z(\col_prog_n[221] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[222].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[222] ),
    .S(write_enable_i),
    .Z(\col_prog_n[222] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[223].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[223] ),
    .S(write_enable_i),
    .Z(\col_prog_n[223] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[224].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[224] ),
    .S(write_enable_i),
    .Z(\col_prog_n[224] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[225].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[225] ),
    .S(write_enable_i),
    .Z(\col_prog_n[225] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[226].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[226] ),
    .S(write_enable_i),
    .Z(\col_prog_n[226] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[227].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[227] ),
    .S(write_enable_i),
    .Z(\col_prog_n[227] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[228].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[228] ),
    .S(write_enable_i),
    .Z(\col_prog_n[228] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[229].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[229] ),
    .S(write_enable_i),
    .Z(\col_prog_n[229] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[22].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[22] ),
    .S(write_enable_i),
    .Z(\col_prog_n[22] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[230].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[230] ),
    .S(write_enable_i),
    .Z(\col_prog_n[230] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[231].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[231] ),
    .S(write_enable_i),
    .Z(\col_prog_n[231] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[232].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[232] ),
    .S(write_enable_i),
    .Z(\col_prog_n[232] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[233].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[233] ),
    .S(write_enable_i),
    .Z(\col_prog_n[233] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[234].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[234] ),
    .S(write_enable_i),
    .Z(\col_prog_n[234] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[235].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[235] ),
    .S(write_enable_i),
    .Z(\col_prog_n[235] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[236].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[236] ),
    .S(write_enable_i),
    .Z(\col_prog_n[236] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[237].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[237] ),
    .S(write_enable_i),
    .Z(\col_prog_n[237] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[238].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[238] ),
    .S(write_enable_i),
    .Z(\col_prog_n[238] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[239].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[239] ),
    .S(write_enable_i),
    .Z(\col_prog_n[239] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[23].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[23] ),
    .S(write_enable_i),
    .Z(\col_prog_n[23] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[240].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[240] ),
    .S(write_enable_i),
    .Z(\col_prog_n[240] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[241].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[241] ),
    .S(write_enable_i),
    .Z(\col_prog_n[241] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[242].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[242] ),
    .S(write_enable_i),
    .Z(\col_prog_n[242] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[243].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[243] ),
    .S(write_enable_i),
    .Z(\col_prog_n[243] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[244].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[244] ),
    .S(write_enable_i),
    .Z(\col_prog_n[244] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[245].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[245] ),
    .S(write_enable_i),
    .Z(\col_prog_n[245] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[246].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[246] ),
    .S(write_enable_i),
    .Z(\col_prog_n[246] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[247].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[247] ),
    .S(write_enable_i),
    .Z(\col_prog_n[247] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[248].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[248] ),
    .S(write_enable_i),
    .Z(\col_prog_n[248] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[249].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[249] ),
    .S(write_enable_i),
    .Z(\col_prog_n[249] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[24].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[24] ),
    .S(write_enable_i),
    .Z(\col_prog_n[24] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[250].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[250] ),
    .S(write_enable_i),
    .Z(\col_prog_n[250] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[251].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[251] ),
    .S(write_enable_i),
    .Z(\col_prog_n[251] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[252].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[252] ),
    .S(write_enable_i),
    .Z(\col_prog_n[252] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[253].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[253] ),
    .S(write_enable_i),
    .Z(\col_prog_n[253] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[254].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[254] ),
    .S(write_enable_i),
    .Z(\col_prog_n[254] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[255].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[255] ),
    .S(write_enable_i),
    .Z(\col_prog_n[255] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[256].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[256] ),
    .S(write_enable_i),
    .Z(\col_prog_n[256] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[257].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[257] ),
    .S(write_enable_i),
    .Z(\col_prog_n[257] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[258].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[258] ),
    .S(write_enable_i),
    .Z(\col_prog_n[258] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[259].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[259] ),
    .S(write_enable_i),
    .Z(\col_prog_n[259] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[25].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[25] ),
    .S(write_enable_i),
    .Z(\col_prog_n[25] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[260].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[260] ),
    .S(write_enable_i),
    .Z(\col_prog_n[260] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[261].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[261] ),
    .S(write_enable_i),
    .Z(\col_prog_n[261] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[262].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[262] ),
    .S(write_enable_i),
    .Z(\col_prog_n[262] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[263].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[263] ),
    .S(write_enable_i),
    .Z(\col_prog_n[263] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[264].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[264] ),
    .S(write_enable_i),
    .Z(\col_prog_n[264] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[265].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[265] ),
    .S(write_enable_i),
    .Z(\col_prog_n[265] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[266].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[266] ),
    .S(write_enable_i),
    .Z(\col_prog_n[266] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[267].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[267] ),
    .S(write_enable_i),
    .Z(\col_prog_n[267] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[268].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[268] ),
    .S(write_enable_i),
    .Z(\col_prog_n[268] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[269].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[269] ),
    .S(write_enable_i),
    .Z(\col_prog_n[269] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[26].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[26] ),
    .S(write_enable_i),
    .Z(\col_prog_n[26] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[270].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[270] ),
    .S(write_enable_i),
    .Z(\col_prog_n[270] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[271].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[271] ),
    .S(write_enable_i),
    .Z(\col_prog_n[271] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[272].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[272] ),
    .S(write_enable_i),
    .Z(\col_prog_n[272] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[273].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[273] ),
    .S(write_enable_i),
    .Z(\col_prog_n[273] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[274].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[274] ),
    .S(write_enable_i),
    .Z(\col_prog_n[274] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[275].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[275] ),
    .S(write_enable_i),
    .Z(\col_prog_n[275] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[276].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[276] ),
    .S(write_enable_i),
    .Z(\col_prog_n[276] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[277].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[277] ),
    .S(write_enable_i),
    .Z(\col_prog_n[277] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[278].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[278] ),
    .S(write_enable_i),
    .Z(\col_prog_n[278] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[279].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[279] ),
    .S(write_enable_i),
    .Z(\col_prog_n[279] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[27].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[27] ),
    .S(write_enable_i),
    .Z(\col_prog_n[27] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[280].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[280] ),
    .S(write_enable_i),
    .Z(\col_prog_n[280] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[281].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[281] ),
    .S(write_enable_i),
    .Z(\col_prog_n[281] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[282].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[282] ),
    .S(write_enable_i),
    .Z(\col_prog_n[282] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[283].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[283] ),
    .S(write_enable_i),
    .Z(\col_prog_n[283] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[284].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[284] ),
    .S(write_enable_i),
    .Z(\col_prog_n[284] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[285].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[285] ),
    .S(write_enable_i),
    .Z(\col_prog_n[285] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[286].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[286] ),
    .S(write_enable_i),
    .Z(\col_prog_n[286] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[287].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[287] ),
    .S(write_enable_i),
    .Z(\col_prog_n[287] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[288].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[288] ),
    .S(write_enable_i),
    .Z(\col_prog_n[288] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[289].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[289] ),
    .S(write_enable_i),
    .Z(\col_prog_n[289] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[28].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[28] ),
    .S(write_enable_i),
    .Z(\col_prog_n[28] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[290].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[290] ),
    .S(write_enable_i),
    .Z(\col_prog_n[290] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[291].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[291] ),
    .S(write_enable_i),
    .Z(\col_prog_n[291] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[292].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[292] ),
    .S(write_enable_i),
    .Z(\col_prog_n[292] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[293].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[293] ),
    .S(write_enable_i),
    .Z(\col_prog_n[293] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[294].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[294] ),
    .S(write_enable_i),
    .Z(\col_prog_n[294] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[295].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[295] ),
    .S(write_enable_i),
    .Z(\col_prog_n[295] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[296].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[296] ),
    .S(write_enable_i),
    .Z(\col_prog_n[296] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[297].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[297] ),
    .S(write_enable_i),
    .Z(\col_prog_n[297] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[298].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[298] ),
    .S(write_enable_i),
    .Z(\col_prog_n[298] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[299].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[299] ),
    .S(write_enable_i),
    .Z(\col_prog_n[299] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[29].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[29] ),
    .S(write_enable_i),
    .Z(\col_prog_n[29] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[2].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[2] ),
    .S(write_enable_i),
    .Z(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[300].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[300] ),
    .S(write_enable_i),
    .Z(\col_prog_n[300] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[301].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[301] ),
    .S(write_enable_i),
    .Z(\col_prog_n[301] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[302].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[302] ),
    .S(write_enable_i),
    .Z(\col_prog_n[302] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[303].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[303] ),
    .S(write_enable_i),
    .Z(\col_prog_n[303] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[304].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[304] ),
    .S(write_enable_i),
    .Z(\col_prog_n[304] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[305].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[305] ),
    .S(write_enable_i),
    .Z(\col_prog_n[305] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[306].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[306] ),
    .S(write_enable_i),
    .Z(\col_prog_n[306] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[307].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[307] ),
    .S(write_enable_i),
    .Z(\col_prog_n[307] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[308].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[308] ),
    .S(write_enable_i),
    .Z(\col_prog_n[308] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[309].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[309] ),
    .S(write_enable_i),
    .Z(\col_prog_n[309] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[30].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[30] ),
    .S(write_enable_i),
    .Z(\col_prog_n[30] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[310].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[310] ),
    .S(write_enable_i),
    .Z(\col_prog_n[310] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[311].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[311] ),
    .S(write_enable_i),
    .Z(\col_prog_n[311] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[312].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[312] ),
    .S(write_enable_i),
    .Z(\col_prog_n[312] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[313].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[313] ),
    .S(write_enable_i),
    .Z(\col_prog_n[313] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[314].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[314] ),
    .S(write_enable_i),
    .Z(\col_prog_n[314] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[315].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[315] ),
    .S(write_enable_i),
    .Z(\col_prog_n[315] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[316].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[316] ),
    .S(write_enable_i),
    .Z(\col_prog_n[316] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[317].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[317] ),
    .S(write_enable_i),
    .Z(\col_prog_n[317] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[318].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[318] ),
    .S(write_enable_i),
    .Z(\col_prog_n[318] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[319].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[319] ),
    .S(write_enable_i),
    .Z(\col_prog_n[319] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[31].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[31] ),
    .S(write_enable_i),
    .Z(\col_prog_n[31] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[320].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[320] ),
    .S(write_enable_i),
    .Z(\col_prog_n[320] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[321].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[321] ),
    .S(write_enable_i),
    .Z(\col_prog_n[321] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[322].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[322] ),
    .S(write_enable_i),
    .Z(\col_prog_n[322] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[323].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[323] ),
    .S(write_enable_i),
    .Z(\col_prog_n[323] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[324].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[324] ),
    .S(write_enable_i),
    .Z(\col_prog_n[324] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[325].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[325] ),
    .S(write_enable_i),
    .Z(\col_prog_n[325] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[326].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[326] ),
    .S(write_enable_i),
    .Z(\col_prog_n[326] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[327].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[327] ),
    .S(write_enable_i),
    .Z(\col_prog_n[327] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[328].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[328] ),
    .S(write_enable_i),
    .Z(\col_prog_n[328] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[329].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[329] ),
    .S(write_enable_i),
    .Z(\col_prog_n[329] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[32].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[32] ),
    .S(write_enable_i),
    .Z(\col_prog_n[32] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[330].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[330] ),
    .S(write_enable_i),
    .Z(\col_prog_n[330] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[331].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[331] ),
    .S(write_enable_i),
    .Z(\col_prog_n[331] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[332].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[332] ),
    .S(write_enable_i),
    .Z(\col_prog_n[332] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[333].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[333] ),
    .S(write_enable_i),
    .Z(\col_prog_n[333] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[334].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[334] ),
    .S(write_enable_i),
    .Z(\col_prog_n[334] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[335].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[335] ),
    .S(write_enable_i),
    .Z(\col_prog_n[335] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[336].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[336] ),
    .S(write_enable_i),
    .Z(\col_prog_n[336] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[337].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[337] ),
    .S(write_enable_i),
    .Z(\col_prog_n[337] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[338].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[338] ),
    .S(write_enable_i),
    .Z(\col_prog_n[338] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[339].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[339] ),
    .S(write_enable_i),
    .Z(\col_prog_n[339] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[33].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[33] ),
    .S(write_enable_i),
    .Z(\col_prog_n[33] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[340].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[340] ),
    .S(write_enable_i),
    .Z(\col_prog_n[340] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[341].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[341] ),
    .S(write_enable_i),
    .Z(\col_prog_n[341] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[342].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[342] ),
    .S(write_enable_i),
    .Z(\col_prog_n[342] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[343].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[343] ),
    .S(write_enable_i),
    .Z(\col_prog_n[343] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[344].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[344] ),
    .S(write_enable_i),
    .Z(\col_prog_n[344] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[345].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[345] ),
    .S(write_enable_i),
    .Z(\col_prog_n[345] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[346].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[346] ),
    .S(write_enable_i),
    .Z(\col_prog_n[346] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[347].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[347] ),
    .S(write_enable_i),
    .Z(\col_prog_n[347] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[348].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[348] ),
    .S(write_enable_i),
    .Z(\col_prog_n[348] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[349].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[349] ),
    .S(write_enable_i),
    .Z(\col_prog_n[349] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[34].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[34] ),
    .S(write_enable_i),
    .Z(\col_prog_n[34] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[350].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[350] ),
    .S(write_enable_i),
    .Z(\col_prog_n[350] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[351].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[351] ),
    .S(write_enable_i),
    .Z(\col_prog_n[351] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[352].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[352] ),
    .S(write_enable_i),
    .Z(\col_prog_n[352] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[353].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[353] ),
    .S(write_enable_i),
    .Z(\col_prog_n[353] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[354].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[354] ),
    .S(write_enable_i),
    .Z(\col_prog_n[354] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[355].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[355] ),
    .S(write_enable_i),
    .Z(\col_prog_n[355] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[356].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[356] ),
    .S(write_enable_i),
    .Z(\col_prog_n[356] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[357].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[357] ),
    .S(write_enable_i),
    .Z(\col_prog_n[357] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[358].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[358] ),
    .S(write_enable_i),
    .Z(\col_prog_n[358] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[359].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[359] ),
    .S(write_enable_i),
    .Z(\col_prog_n[359] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[35].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[35] ),
    .S(write_enable_i),
    .Z(\col_prog_n[35] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[360].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[360] ),
    .S(write_enable_i),
    .Z(\col_prog_n[360] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[361].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[361] ),
    .S(write_enable_i),
    .Z(\col_prog_n[361] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[362].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[362] ),
    .S(write_enable_i),
    .Z(\col_prog_n[362] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[363].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[363] ),
    .S(write_enable_i),
    .Z(\col_prog_n[363] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[364].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[364] ),
    .S(write_enable_i),
    .Z(\col_prog_n[364] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[365].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[365] ),
    .S(write_enable_i),
    .Z(\col_prog_n[365] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[366].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[366] ),
    .S(write_enable_i),
    .Z(\col_prog_n[366] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[367].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[367] ),
    .S(write_enable_i),
    .Z(\col_prog_n[367] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[368].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[368] ),
    .S(write_enable_i),
    .Z(\col_prog_n[368] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[369].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[369] ),
    .S(write_enable_i),
    .Z(\col_prog_n[369] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[36].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[36] ),
    .S(write_enable_i),
    .Z(\col_prog_n[36] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[370].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[370] ),
    .S(write_enable_i),
    .Z(\col_prog_n[370] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[371].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[371] ),
    .S(write_enable_i),
    .Z(\col_prog_n[371] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[372].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[372] ),
    .S(write_enable_i),
    .Z(\col_prog_n[372] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[373].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[373] ),
    .S(write_enable_i),
    .Z(\col_prog_n[373] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[374].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[374] ),
    .S(write_enable_i),
    .Z(\col_prog_n[374] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[375].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[375] ),
    .S(write_enable_i),
    .Z(\col_prog_n[375] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[376].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[376] ),
    .S(write_enable_i),
    .Z(\col_prog_n[376] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[377].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[377] ),
    .S(write_enable_i),
    .Z(\col_prog_n[377] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[378].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[378] ),
    .S(write_enable_i),
    .Z(\col_prog_n[378] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[379].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[379] ),
    .S(write_enable_i),
    .Z(\col_prog_n[379] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[37].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[37] ),
    .S(write_enable_i),
    .Z(\col_prog_n[37] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[380].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[380] ),
    .S(write_enable_i),
    .Z(\col_prog_n[380] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[381].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[381] ),
    .S(write_enable_i),
    .Z(\col_prog_n[381] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[382].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[382] ),
    .S(write_enable_i),
    .Z(\col_prog_n[382] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[383].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[383] ),
    .S(write_enable_i),
    .Z(\col_prog_n[383] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[384].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[384] ),
    .S(write_enable_i),
    .Z(\col_prog_n[384] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[385].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[385] ),
    .S(write_enable_i),
    .Z(\col_prog_n[385] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[386].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[386] ),
    .S(write_enable_i),
    .Z(\col_prog_n[386] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[387].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[387] ),
    .S(write_enable_i),
    .Z(\col_prog_n[387] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[388].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[388] ),
    .S(write_enable_i),
    .Z(\col_prog_n[388] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[389].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[389] ),
    .S(write_enable_i),
    .Z(\col_prog_n[389] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[38].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[38] ),
    .S(write_enable_i),
    .Z(\col_prog_n[38] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[390].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[390] ),
    .S(write_enable_i),
    .Z(\col_prog_n[390] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[391].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[391] ),
    .S(write_enable_i),
    .Z(\col_prog_n[391] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[392].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[392] ),
    .S(write_enable_i),
    .Z(\col_prog_n[392] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[393].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[393] ),
    .S(write_enable_i),
    .Z(\col_prog_n[393] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[394].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[394] ),
    .S(write_enable_i),
    .Z(\col_prog_n[394] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[395].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[395] ),
    .S(write_enable_i),
    .Z(\col_prog_n[395] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[396].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[396] ),
    .S(write_enable_i),
    .Z(\col_prog_n[396] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[397].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[397] ),
    .S(write_enable_i),
    .Z(\col_prog_n[397] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[398].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[398] ),
    .S(write_enable_i),
    .Z(\col_prog_n[398] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[399].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[399] ),
    .S(write_enable_i),
    .Z(\col_prog_n[399] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[39].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[39] ),
    .S(write_enable_i),
    .Z(\col_prog_n[39] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[3].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[3] ),
    .S(write_enable_i),
    .Z(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[400].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[400] ),
    .S(write_enable_i),
    .Z(\col_prog_n[400] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[401].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[401] ),
    .S(write_enable_i),
    .Z(\col_prog_n[401] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[402].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[402] ),
    .S(write_enable_i),
    .Z(\col_prog_n[402] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[403].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[403] ),
    .S(write_enable_i),
    .Z(\col_prog_n[403] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[404].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[404] ),
    .S(write_enable_i),
    .Z(\col_prog_n[404] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[405].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[405] ),
    .S(write_enable_i),
    .Z(\col_prog_n[405] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[406].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[406] ),
    .S(write_enable_i),
    .Z(\col_prog_n[406] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[407].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[407] ),
    .S(write_enable_i),
    .Z(\col_prog_n[407] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[408].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[408] ),
    .S(write_enable_i),
    .Z(\col_prog_n[408] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[409].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[409] ),
    .S(write_enable_i),
    .Z(\col_prog_n[409] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[40].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[40] ),
    .S(write_enable_i),
    .Z(\col_prog_n[40] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[410].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[410] ),
    .S(write_enable_i),
    .Z(\col_prog_n[410] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[411].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[411] ),
    .S(write_enable_i),
    .Z(\col_prog_n[411] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[412].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[412] ),
    .S(write_enable_i),
    .Z(\col_prog_n[412] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[413].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[413] ),
    .S(write_enable_i),
    .Z(\col_prog_n[413] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[414].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[414] ),
    .S(write_enable_i),
    .Z(\col_prog_n[414] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[415].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[415] ),
    .S(write_enable_i),
    .Z(\col_prog_n[415] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[416].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[416] ),
    .S(write_enable_i),
    .Z(\col_prog_n[416] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[417].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[417] ),
    .S(write_enable_i),
    .Z(\col_prog_n[417] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[418].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[418] ),
    .S(write_enable_i),
    .Z(\col_prog_n[418] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[419].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[419] ),
    .S(write_enable_i),
    .Z(\col_prog_n[419] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[41].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[41] ),
    .S(write_enable_i),
    .Z(\col_prog_n[41] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[420].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[420] ),
    .S(write_enable_i),
    .Z(\col_prog_n[420] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[421].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[421] ),
    .S(write_enable_i),
    .Z(\col_prog_n[421] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[422].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[422] ),
    .S(write_enable_i),
    .Z(\col_prog_n[422] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[423].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[423] ),
    .S(write_enable_i),
    .Z(\col_prog_n[423] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[424].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[424] ),
    .S(write_enable_i),
    .Z(\col_prog_n[424] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[425].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[425] ),
    .S(write_enable_i),
    .Z(\col_prog_n[425] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[426].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[426] ),
    .S(write_enable_i),
    .Z(\col_prog_n[426] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[427].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[427] ),
    .S(write_enable_i),
    .Z(\col_prog_n[427] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[428].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[428] ),
    .S(write_enable_i),
    .Z(\col_prog_n[428] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[429].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[429] ),
    .S(write_enable_i),
    .Z(\col_prog_n[429] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[42].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[42] ),
    .S(write_enable_i),
    .Z(\col_prog_n[42] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[430].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[430] ),
    .S(write_enable_i),
    .Z(\col_prog_n[430] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[431].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[431] ),
    .S(write_enable_i),
    .Z(\col_prog_n[431] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[432].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[432] ),
    .S(write_enable_i),
    .Z(\col_prog_n[432] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[433].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[433] ),
    .S(write_enable_i),
    .Z(\col_prog_n[433] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[434].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[434] ),
    .S(write_enable_i),
    .Z(\col_prog_n[434] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[435].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[435] ),
    .S(write_enable_i),
    .Z(\col_prog_n[435] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[436].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[436] ),
    .S(write_enable_i),
    .Z(\col_prog_n[436] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[437].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[437] ),
    .S(write_enable_i),
    .Z(\col_prog_n[437] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[438].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[438] ),
    .S(write_enable_i),
    .Z(\col_prog_n[438] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[439].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[439] ),
    .S(write_enable_i),
    .Z(\col_prog_n[439] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[43].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[43] ),
    .S(write_enable_i),
    .Z(\col_prog_n[43] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[440].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[440] ),
    .S(write_enable_i),
    .Z(\col_prog_n[440] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[441].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[441] ),
    .S(write_enable_i),
    .Z(\col_prog_n[441] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[442].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[442] ),
    .S(write_enable_i),
    .Z(\col_prog_n[442] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[443].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[443] ),
    .S(write_enable_i),
    .Z(\col_prog_n[443] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[444].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[444] ),
    .S(write_enable_i),
    .Z(\col_prog_n[444] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[445].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[445] ),
    .S(write_enable_i),
    .Z(\col_prog_n[445] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[446].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[446] ),
    .S(write_enable_i),
    .Z(\col_prog_n[446] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[447].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[447] ),
    .S(write_enable_i),
    .Z(\col_prog_n[447] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[448].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[448] ),
    .S(write_enable_i),
    .Z(\col_prog_n[448] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[449].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[449] ),
    .S(write_enable_i),
    .Z(\col_prog_n[449] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[44].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[44] ),
    .S(write_enable_i),
    .Z(\col_prog_n[44] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[450].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[450] ),
    .S(write_enable_i),
    .Z(\col_prog_n[450] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[451].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[451] ),
    .S(write_enable_i),
    .Z(\col_prog_n[451] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[452].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[452] ),
    .S(write_enable_i),
    .Z(\col_prog_n[452] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[453].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[453] ),
    .S(write_enable_i),
    .Z(\col_prog_n[453] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[454].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[454] ),
    .S(write_enable_i),
    .Z(\col_prog_n[454] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[455].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[455] ),
    .S(write_enable_i),
    .Z(\col_prog_n[455] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[456].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[456] ),
    .S(write_enable_i),
    .Z(\col_prog_n[456] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[457].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[457] ),
    .S(write_enable_i),
    .Z(\col_prog_n[457] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[458].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[458] ),
    .S(write_enable_i),
    .Z(\col_prog_n[458] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[459].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[459] ),
    .S(write_enable_i),
    .Z(\col_prog_n[459] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[45].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[45] ),
    .S(write_enable_i),
    .Z(\col_prog_n[45] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[460].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[460] ),
    .S(write_enable_i),
    .Z(\col_prog_n[460] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[461].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[461] ),
    .S(write_enable_i),
    .Z(\col_prog_n[461] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[462].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[462] ),
    .S(write_enable_i),
    .Z(\col_prog_n[462] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[463].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[463] ),
    .S(write_enable_i),
    .Z(\col_prog_n[463] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[464].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[464] ),
    .S(write_enable_i),
    .Z(\col_prog_n[464] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[465].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[465] ),
    .S(write_enable_i),
    .Z(\col_prog_n[465] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[466].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[466] ),
    .S(write_enable_i),
    .Z(\col_prog_n[466] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[467].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[467] ),
    .S(write_enable_i),
    .Z(\col_prog_n[467] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[468].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[468] ),
    .S(write_enable_i),
    .Z(\col_prog_n[468] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[469].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[469] ),
    .S(write_enable_i),
    .Z(\col_prog_n[469] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[46].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[46] ),
    .S(write_enable_i),
    .Z(\col_prog_n[46] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[470].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[470] ),
    .S(write_enable_i),
    .Z(\col_prog_n[470] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[471].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[471] ),
    .S(write_enable_i),
    .Z(\col_prog_n[471] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[472].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[472] ),
    .S(write_enable_i),
    .Z(\col_prog_n[472] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[473].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[473] ),
    .S(write_enable_i),
    .Z(\col_prog_n[473] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[474].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[474] ),
    .S(write_enable_i),
    .Z(\col_prog_n[474] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[475].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[475] ),
    .S(write_enable_i),
    .Z(\col_prog_n[475] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[476].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[476] ),
    .S(write_enable_i),
    .Z(\col_prog_n[476] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[477].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[477] ),
    .S(write_enable_i),
    .Z(\col_prog_n[477] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[478].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[478] ),
    .S(write_enable_i),
    .Z(\col_prog_n[478] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[479].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[479] ),
    .S(write_enable_i),
    .Z(\col_prog_n[479] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[47].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[47] ),
    .S(write_enable_i),
    .Z(\col_prog_n[47] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[480].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[480] ),
    .S(write_enable_i),
    .Z(\col_prog_n[480] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[481].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[481] ),
    .S(write_enable_i),
    .Z(\col_prog_n[481] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[482].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[482] ),
    .S(write_enable_i),
    .Z(\col_prog_n[482] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[483].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[483] ),
    .S(write_enable_i),
    .Z(\col_prog_n[483] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[484].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[484] ),
    .S(write_enable_i),
    .Z(\col_prog_n[484] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[485].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[485] ),
    .S(write_enable_i),
    .Z(\col_prog_n[485] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[486].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[486] ),
    .S(write_enable_i),
    .Z(\col_prog_n[486] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[487].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[487] ),
    .S(write_enable_i),
    .Z(\col_prog_n[487] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[488].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[488] ),
    .S(write_enable_i),
    .Z(\col_prog_n[488] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[489].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[489] ),
    .S(write_enable_i),
    .Z(\col_prog_n[489] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[48].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[48] ),
    .S(write_enable_i),
    .Z(\col_prog_n[48] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[490].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[490] ),
    .S(write_enable_i),
    .Z(\col_prog_n[490] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[491].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[491] ),
    .S(write_enable_i),
    .Z(\col_prog_n[491] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[492].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[492] ),
    .S(write_enable_i),
    .Z(\col_prog_n[492] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[493].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[493] ),
    .S(write_enable_i),
    .Z(\col_prog_n[493] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[494].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[494] ),
    .S(write_enable_i),
    .Z(\col_prog_n[494] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[495].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[495] ),
    .S(write_enable_i),
    .Z(\col_prog_n[495] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[496].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[496] ),
    .S(write_enable_i),
    .Z(\col_prog_n[496] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[497].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[497] ),
    .S(write_enable_i),
    .Z(\col_prog_n[497] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[498].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[498] ),
    .S(write_enable_i),
    .Z(\col_prog_n[498] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[499].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[499] ),
    .S(write_enable_i),
    .Z(\col_prog_n[499] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[49].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[49] ),
    .S(write_enable_i),
    .Z(\col_prog_n[49] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[4].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[4] ),
    .S(write_enable_i),
    .Z(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[500].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[500] ),
    .S(write_enable_i),
    .Z(\col_prog_n[500] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[501].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[501] ),
    .S(write_enable_i),
    .Z(\col_prog_n[501] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[502].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[502] ),
    .S(write_enable_i),
    .Z(\col_prog_n[502] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[503].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[503] ),
    .S(write_enable_i),
    .Z(\col_prog_n[503] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[504].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[504] ),
    .S(write_enable_i),
    .Z(\col_prog_n[504] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[505].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[505] ),
    .S(write_enable_i),
    .Z(\col_prog_n[505] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[506].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[506] ),
    .S(write_enable_i),
    .Z(\col_prog_n[506] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[507].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[507] ),
    .S(write_enable_i),
    .Z(\col_prog_n[507] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[508].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[508] ),
    .S(write_enable_i),
    .Z(\col_prog_n[508] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[509].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[509] ),
    .S(write_enable_i),
    .Z(\col_prog_n[509] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[50].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[50] ),
    .S(write_enable_i),
    .Z(\col_prog_n[50] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[510].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[510] ),
    .S(write_enable_i),
    .Z(\col_prog_n[510] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[511].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[511] ),
    .S(write_enable_i),
    .Z(\col_prog_n[511] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[51].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[51] ),
    .S(write_enable_i),
    .Z(\col_prog_n[51] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[52].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[52] ),
    .S(write_enable_i),
    .Z(\col_prog_n[52] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[53].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[53] ),
    .S(write_enable_i),
    .Z(\col_prog_n[53] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[54].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[54] ),
    .S(write_enable_i),
    .Z(\col_prog_n[54] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[55].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[55] ),
    .S(write_enable_i),
    .Z(\col_prog_n[55] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[56].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[56] ),
    .S(write_enable_i),
    .Z(\col_prog_n[56] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[57].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[57] ),
    .S(write_enable_i),
    .Z(\col_prog_n[57] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[58].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[58] ),
    .S(write_enable_i),
    .Z(\col_prog_n[58] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[59].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[59] ),
    .S(write_enable_i),
    .Z(\col_prog_n[59] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[5].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[5] ),
    .S(write_enable_i),
    .Z(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[60].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[60] ),
    .S(write_enable_i),
    .Z(\col_prog_n[60] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[61].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[61] ),
    .S(write_enable_i),
    .Z(\col_prog_n[61] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[62].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[62] ),
    .S(write_enable_i),
    .Z(\col_prog_n[62] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[63].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[63] ),
    .S(write_enable_i),
    .Z(\col_prog_n[63] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[64].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[64] ),
    .S(write_enable_i),
    .Z(\col_prog_n[64] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[65].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[65] ),
    .S(write_enable_i),
    .Z(\col_prog_n[65] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[66].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[66] ),
    .S(write_enable_i),
    .Z(\col_prog_n[66] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[67].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[67] ),
    .S(write_enable_i),
    .Z(\col_prog_n[67] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[68].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[68] ),
    .S(write_enable_i),
    .Z(\col_prog_n[68] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[69].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[69] ),
    .S(write_enable_i),
    .Z(\col_prog_n[69] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[6].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[6] ),
    .S(write_enable_i),
    .Z(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[70].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[70] ),
    .S(write_enable_i),
    .Z(\col_prog_n[70] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[71].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[71] ),
    .S(write_enable_i),
    .Z(\col_prog_n[71] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[72].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[72] ),
    .S(write_enable_i),
    .Z(\col_prog_n[72] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[73].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[73] ),
    .S(write_enable_i),
    .Z(\col_prog_n[73] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[74].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[74] ),
    .S(write_enable_i),
    .Z(\col_prog_n[74] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[75].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[75] ),
    .S(write_enable_i),
    .Z(\col_prog_n[75] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[76].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[76] ),
    .S(write_enable_i),
    .Z(\col_prog_n[76] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[77].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[77] ),
    .S(write_enable_i),
    .Z(\col_prog_n[77] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[78].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[78] ),
    .S(write_enable_i),
    .Z(\col_prog_n[78] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[79].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[79] ),
    .S(write_enable_i),
    .Z(\col_prog_n[79] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[7].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[7] ),
    .S(write_enable_i),
    .Z(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[80].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[80] ),
    .S(write_enable_i),
    .Z(\col_prog_n[80] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[81].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[81] ),
    .S(write_enable_i),
    .Z(\col_prog_n[81] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[82].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[82] ),
    .S(write_enable_i),
    .Z(\col_prog_n[82] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[83].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[83] ),
    .S(write_enable_i),
    .Z(\col_prog_n[83] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[84].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[84] ),
    .S(write_enable_i),
    .Z(\col_prog_n[84] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[85].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[85] ),
    .S(write_enable_i),
    .Z(\col_prog_n[85] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[86].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[86] ),
    .S(write_enable_i),
    .Z(\col_prog_n[86] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[87].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[87] ),
    .S(write_enable_i),
    .Z(\col_prog_n[87] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[88].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[88] ),
    .S(write_enable_i),
    .Z(\col_prog_n[88] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[89].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[89] ),
    .S(write_enable_i),
    .Z(\col_prog_n[89] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[8].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[8] ),
    .S(write_enable_i),
    .Z(\col_prog_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[90].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[90] ),
    .S(write_enable_i),
    .Z(\col_prog_n[90] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[91].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[91] ),
    .S(write_enable_i),
    .Z(\col_prog_n[91] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[92].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[92] ),
    .S(write_enable_i),
    .Z(\col_prog_n[92] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[93].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[93] ),
    .S(write_enable_i),
    .Z(\col_prog_n[93] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[94].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[94] ),
    .S(write_enable_i),
    .Z(\col_prog_n[94] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[95].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[95] ),
    .S(write_enable_i),
    .Z(\col_prog_n[95] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[96].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[96] ),
    .S(write_enable_i),
    .Z(\col_prog_n[96] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[97].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[97] ),
    .S(write_enable_i),
    .Z(\col_prog_n[97] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[98].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[98] ),
    .S(write_enable_i),
    .Z(\col_prog_n[98] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[99].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[99] ),
    .S(write_enable_i),
    .Z(\col_prog_n[99] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 \genblk2[9].prog_disable_keep_cell  (.I0(one),
    .I1(\col_prog_n_reg[9] ),
    .S(write_enable_i),
    .Z(\col_prog_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[0].bitsel_buf_keep_cell  (.I(\bit_sel_reg[0] ),
    .Z(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[10].bitsel_buf_keep_cell  (.I(\bit_sel_reg[10] ),
    .Z(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[11].bitsel_buf_keep_cell  (.I(\bit_sel_reg[11] ),
    .Z(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[12].bitsel_buf_keep_cell  (.I(\bit_sel_reg[12] ),
    .Z(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[13].bitsel_buf_keep_cell  (.I(\bit_sel_reg[13] ),
    .Z(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[14].bitsel_buf_keep_cell  (.I(\bit_sel_reg[14] ),
    .Z(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[15].bitsel_buf_keep_cell  (.I(\bit_sel_reg[15] ),
    .Z(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[16].bitsel_buf_keep_cell  (.I(\bit_sel_reg[16] ),
    .Z(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[17].bitsel_buf_keep_cell  (.I(\bit_sel_reg[17] ),
    .Z(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[18].bitsel_buf_keep_cell  (.I(\bit_sel_reg[18] ),
    .Z(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[19].bitsel_buf_keep_cell  (.I(\bit_sel_reg[19] ),
    .Z(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[1].bitsel_buf_keep_cell  (.I(\bit_sel_reg[1] ),
    .Z(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[20].bitsel_buf_keep_cell  (.I(\bit_sel_reg[20] ),
    .Z(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[21].bitsel_buf_keep_cell  (.I(\bit_sel_reg[21] ),
    .Z(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[22].bitsel_buf_keep_cell  (.I(\bit_sel_reg[22] ),
    .Z(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[23].bitsel_buf_keep_cell  (.I(\bit_sel_reg[23] ),
    .Z(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[24].bitsel_buf_keep_cell  (.I(\bit_sel_reg[24] ),
    .Z(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[25].bitsel_buf_keep_cell  (.I(\bit_sel_reg[25] ),
    .Z(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[26].bitsel_buf_keep_cell  (.I(\bit_sel_reg[26] ),
    .Z(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[27].bitsel_buf_keep_cell  (.I(\bit_sel_reg[27] ),
    .Z(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[28].bitsel_buf_keep_cell  (.I(\bit_sel_reg[28] ),
    .Z(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[29].bitsel_buf_keep_cell  (.I(\bit_sel_reg[29] ),
    .Z(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[2].bitsel_buf_keep_cell  (.I(\bit_sel_reg[2] ),
    .Z(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[30].bitsel_buf_keep_cell  (.I(\bit_sel_reg[30] ),
    .Z(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[31].bitsel_buf_keep_cell  (.I(\bit_sel_reg[31] ),
    .Z(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[32].bitsel_buf_keep_cell  (.I(\bit_sel_reg[32] ),
    .Z(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[33].bitsel_buf_keep_cell  (.I(\bit_sel_reg[33] ),
    .Z(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[34].bitsel_buf_keep_cell  (.I(\bit_sel_reg[34] ),
    .Z(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[35].bitsel_buf_keep_cell  (.I(\bit_sel_reg[35] ),
    .Z(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[36].bitsel_buf_keep_cell  (.I(\bit_sel_reg[36] ),
    .Z(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[37].bitsel_buf_keep_cell  (.I(\bit_sel_reg[37] ),
    .Z(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[38].bitsel_buf_keep_cell  (.I(\bit_sel_reg[38] ),
    .Z(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[39].bitsel_buf_keep_cell  (.I(\bit_sel_reg[39] ),
    .Z(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[3].bitsel_buf_keep_cell  (.I(\bit_sel_reg[3] ),
    .Z(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[40].bitsel_buf_keep_cell  (.I(\bit_sel_reg[40] ),
    .Z(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[41].bitsel_buf_keep_cell  (.I(\bit_sel_reg[41] ),
    .Z(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[42].bitsel_buf_keep_cell  (.I(\bit_sel_reg[42] ),
    .Z(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[43].bitsel_buf_keep_cell  (.I(\bit_sel_reg[43] ),
    .Z(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[44].bitsel_buf_keep_cell  (.I(\bit_sel_reg[44] ),
    .Z(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[45].bitsel_buf_keep_cell  (.I(\bit_sel_reg[45] ),
    .Z(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[46].bitsel_buf_keep_cell  (.I(\bit_sel_reg[46] ),
    .Z(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[47].bitsel_buf_keep_cell  (.I(\bit_sel_reg[47] ),
    .Z(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[48].bitsel_buf_keep_cell  (.I(\bit_sel_reg[48] ),
    .Z(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[49].bitsel_buf_keep_cell  (.I(\bit_sel_reg[49] ),
    .Z(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[4].bitsel_buf_keep_cell  (.I(\bit_sel_reg[4] ),
    .Z(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[50].bitsel_buf_keep_cell  (.I(\bit_sel_reg[50] ),
    .Z(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[51].bitsel_buf_keep_cell  (.I(\bit_sel_reg[51] ),
    .Z(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[52].bitsel_buf_keep_cell  (.I(\bit_sel_reg[52] ),
    .Z(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[53].bitsel_buf_keep_cell  (.I(\bit_sel_reg[53] ),
    .Z(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[54].bitsel_buf_keep_cell  (.I(\bit_sel_reg[54] ),
    .Z(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[55].bitsel_buf_keep_cell  (.I(\bit_sel_reg[55] ),
    .Z(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[56].bitsel_buf_keep_cell  (.I(\bit_sel_reg[56] ),
    .Z(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[57].bitsel_buf_keep_cell  (.I(\bit_sel_reg[57] ),
    .Z(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[58].bitsel_buf_keep_cell  (.I(\bit_sel_reg[58] ),
    .Z(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[59].bitsel_buf_keep_cell  (.I(\bit_sel_reg[59] ),
    .Z(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[5].bitsel_buf_keep_cell  (.I(\bit_sel_reg[5] ),
    .Z(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[60].bitsel_buf_keep_cell  (.I(\bit_sel_reg[60] ),
    .Z(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[61].bitsel_buf_keep_cell  (.I(\bit_sel_reg[61] ),
    .Z(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[62].bitsel_buf_keep_cell  (.I(\bit_sel_reg[62] ),
    .Z(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[63].bitsel_buf_keep_cell  (.I(\bit_sel_reg[63] ),
    .Z(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[6].bitsel_buf_keep_cell  (.I(\bit_sel_reg[6] ),
    .Z(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[7].bitsel_buf_keep_cell  (.I(\bit_sel_reg[7] ),
    .Z(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[8].bitsel_buf_keep_cell  (.I(\bit_sel_reg[8] ),
    .Z(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk3[9].bitsel_buf_keep_cell  (.I(\bit_sel_reg[9] ),
    .Z(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].preset_buf_keep_cell  (.I(\preset_n_reg[0] ),
    .Z(\preset_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[0].sense_buf_keep_cell  (.I(\sense_del[0] ),
    .Z(\sense[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[0].sense_dly_keep_cell  (.I(\sense_reg[0] ),
    .Z(\sense_del[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[10].preset_buf_keep_cell  (.I(\preset_n_reg[10] ),
    .Z(\preset_n[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[10].sense_buf_keep_cell  (.I(\sense_del[10] ),
    .Z(\sense[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[10].sense_dly_keep_cell  (.I(\sense_reg[10] ),
    .Z(\sense_del[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[11].preset_buf_keep_cell  (.I(\preset_n_reg[11] ),
    .Z(\preset_n[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[11].sense_buf_keep_cell  (.I(\sense_del[11] ),
    .Z(\sense[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[11].sense_dly_keep_cell  (.I(\sense_reg[11] ),
    .Z(\sense_del[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[12].preset_buf_keep_cell  (.I(\preset_n_reg[12] ),
    .Z(\preset_n[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[12].sense_buf_keep_cell  (.I(\sense_del[12] ),
    .Z(\sense[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[12].sense_dly_keep_cell  (.I(\sense_reg[12] ),
    .Z(\sense_del[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[13].preset_buf_keep_cell  (.I(\preset_n_reg[13] ),
    .Z(\preset_n[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[13].sense_buf_keep_cell  (.I(\sense_del[13] ),
    .Z(\sense[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[13].sense_dly_keep_cell  (.I(\sense_reg[13] ),
    .Z(\sense_del[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[14].preset_buf_keep_cell  (.I(\preset_n_reg[14] ),
    .Z(\preset_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[14].sense_buf_keep_cell  (.I(\sense_del[14] ),
    .Z(\sense[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[14].sense_dly_keep_cell  (.I(\sense_reg[14] ),
    .Z(\sense_del[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[15].preset_buf_keep_cell  (.I(\preset_n_reg[15] ),
    .Z(\preset_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[15].sense_buf_keep_cell  (.I(\sense_del[15] ),
    .Z(\sense[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[15].sense_dly_keep_cell  (.I(\sense_reg[15] ),
    .Z(\sense_del[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[1].preset_buf_keep_cell  (.I(\preset_n_reg[1] ),
    .Z(\preset_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[1].sense_buf_keep_cell  (.I(\sense_del[1] ),
    .Z(\sense[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[1].sense_dly_keep_cell  (.I(\sense_reg[1] ),
    .Z(\sense_del[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[2].preset_buf_keep_cell  (.I(\preset_n_reg[2] ),
    .Z(\preset_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[2].sense_buf_keep_cell  (.I(\sense_del[2] ),
    .Z(\sense[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[2].sense_dly_keep_cell  (.I(\sense_reg[2] ),
    .Z(\sense_del[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[3].preset_buf_keep_cell  (.I(\preset_n_reg[3] ),
    .Z(\preset_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[3].sense_buf_keep_cell  (.I(\sense_del[3] ),
    .Z(\sense[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[3].sense_dly_keep_cell  (.I(\sense_reg[3] ),
    .Z(\sense_del[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[4].preset_buf_keep_cell  (.I(\preset_n_reg[4] ),
    .Z(\preset_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[4].sense_buf_keep_cell  (.I(\sense_del[4] ),
    .Z(\sense[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[4].sense_dly_keep_cell  (.I(\sense_reg[4] ),
    .Z(\sense_del[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[5].preset_buf_keep_cell  (.I(\preset_n_reg[5] ),
    .Z(\preset_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[5].sense_buf_keep_cell  (.I(\sense_del[5] ),
    .Z(\sense[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[5].sense_dly_keep_cell  (.I(\sense_reg[5] ),
    .Z(\sense_del[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[6].preset_buf_keep_cell  (.I(\preset_n_reg[6] ),
    .Z(\preset_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[6].sense_buf_keep_cell  (.I(\sense_del[6] ),
    .Z(\sense[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[6].sense_dly_keep_cell  (.I(\sense_reg[6] ),
    .Z(\sense_del[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[7].preset_buf_keep_cell  (.I(\preset_n_reg[7] ),
    .Z(\preset_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[7].sense_buf_keep_cell  (.I(\sense_del[7] ),
    .Z(\sense[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[7].sense_dly_keep_cell  (.I(\sense_reg[7] ),
    .Z(\sense_del[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[8].preset_buf_keep_cell  (.I(\preset_n_reg[8] ),
    .Z(\preset_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[8].sense_buf_keep_cell  (.I(\sense_del[8] ),
    .Z(\sense[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[8].sense_dly_keep_cell  (.I(\sense_reg[8] ),
    .Z(\sense_del[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[9].preset_buf_keep_cell  (.I(\preset_n_reg[9] ),
    .Z(\preset_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 \genblk4[9].sense_buf_keep_cell  (.I(\sense_del[9] ),
    .Z(\sense[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_2 \genblk4[9].sense_dly_keep_cell  (.I(\sense_reg[9] ),
    .Z(\sense_del[9] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh tie_keep_cell (.Z(one));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Left_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Left_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Left_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Left_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Left_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Left_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Left_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Left_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Left_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Left_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Left_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Left_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Left_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Left_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Left_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Left_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_2_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_2_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_2_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_2_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_2_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_2_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_2_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_2_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_2_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_2_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_2_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_2_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_2_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_2_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_2_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_2_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_2_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_2_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_2_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_2_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_2_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_2_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_2_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_2_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_2_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_2_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_2_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_2_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_2_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_2_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_2_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_2_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_2_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_2_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_2_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_2_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_2_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_2_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_2_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_2_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_2_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_2_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_2_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_2_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_2_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_2_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_2_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_2_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_2_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_2_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_2_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_2_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_2_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_2_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_2_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_2_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_2_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_2_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_2_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_2_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_2_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_2_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_2_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_2_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_2_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_2_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_2_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_2_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_2_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_2_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_2_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_2_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_2_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_2_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_2_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_2_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_2_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_2_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_2_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_2_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_2_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_2_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_2_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_2_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_2_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_2_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_2_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_2_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_2_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_2_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_2_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_2_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_2_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_2_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_2_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_2_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_2_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_2_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_2_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_2_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_2_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_2_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_2_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_2_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_2_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_2_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_2_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_2_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_2_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_2_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_2_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_2_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_2_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_2_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_2_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_2_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_2_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_2_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_2_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_2_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_2_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_2_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_2_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_2_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_2_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_2_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_2_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_2_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_2_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_2_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_2_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_2_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_2_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_2_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_2_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_2_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_2_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_2_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_2_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_2_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_2_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_2_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_2_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Right_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Right_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Right_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Right_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Right_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Right_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Right_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Right_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Right_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Right_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Right_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Right_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Right_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Right_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Right_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Right_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Right_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Right_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Right_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Right_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Right_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Right_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Right_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Right_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Right_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Right_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Right_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Right_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Right_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Right_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Right_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Right_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Right_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Right_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Right_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Right_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Right_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Right_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Right_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Right_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Right_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Right_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Right_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Right_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Right_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Right_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Right_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Right_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Right_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Right_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Right_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Right_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Right_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Right_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Right_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Right_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Right_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Right_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Right_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Right_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Right_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Right_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Right_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Right_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Right_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Right_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Right_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Right_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Right_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Right_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Right_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Right_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Right_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Right_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Right_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Right_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Right_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Right_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Right_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Right_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Right_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Right_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Right_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Right_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Right_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Right_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Right_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Right_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Right_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Right_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Right_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Right_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Right_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Right_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Right_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Right_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Right_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Right_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Right_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Right_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Right_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Right_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Right_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Right_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Right_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Right_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Right_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Right_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Right_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Right_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Right_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Right_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Right_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Right_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Right_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_2_Right_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_2_Right_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_2_Right_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_2_Right_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_2_Right_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_2_Right_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_2_Right_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_2_Right_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_2_Right_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_2_Right_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_2_Right_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_2_Right_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_2_Right_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_2_Right_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_2_Right_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_2_Right_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_2_Right_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_2_Right_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_2_Right_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_2_Right_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_2_Right_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_2_Right_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_2_Right_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_2_Right_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_2_Right_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_2_Right_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_2_Right_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_2_Right_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_2_Right_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_2_Right_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_2_Right_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_2_Right_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_2_Right_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_2_Right_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_2_Right_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_2_Right_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_2_Right_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_2_Right_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_2_Right_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_2_Right_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_2_Right_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_2_Right_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_2_Right_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_2_Right_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_2_Right_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_2_Right_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_2_Right_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_2_Right_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_2_Right_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_2_Right_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_2_Right_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_2_Right_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_2_Right_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_2_Right_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_2_Right_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_2_Right_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_2_Right_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_2_Right_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_2_Right_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_2_Right_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_2_Right_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_2_Right_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_2_Right_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_2_Right_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_2_Right_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_2_Right_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_2_Right_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_2_Right_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_2_Right_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_2_Right_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_2_Right_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_2_Right_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_2_Right_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_2_Right_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_2_Right_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_2_Right_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_2_Right_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_2_Right_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_2_Right_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_2_Right_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_2_Right_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_2_Right_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_2_Right_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_2_Right_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_2_Right_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_2_Right_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_2_Right_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_2_Right_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_2_Right_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_2_Right_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_2_Right_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_2_Right_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_2_Right_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_2_Right_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_2_Right_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_2_Right_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_2_Right_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_2_Right_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_2_Right_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_2_Right_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_2_Right_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_2_Right_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_2_Right_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_2_Right_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_2_Right_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_2_Right_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_2_Right_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_2_Right_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_2_Right_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_2_Right_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_2_Right_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_2_Right_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_2_Right_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_2_Right_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_2_Right_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_2_Right_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_2_Right_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_2_Right_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_2_Right_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_2_Right_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_2_Right_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_2_Right_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_2_Right_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_2_Right_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_2_Right_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_2_Right_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_2_Right_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_2_Right_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_2_Right_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_2_Right_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_2_Right_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_2_Right_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_2_Right_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_2_Right_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_2_Right_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_2_Right_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_2_Right_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_2_Right_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_2_Right_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_2_Right_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_2_Right_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_2_Right_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_2_Right_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Right_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_3_Left_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_3_Left_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_3_Left_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_3_Left_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_3_Left_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_3_Left_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_3_Left_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_3_Left_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_3_Left_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_3_Left_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_3_Left_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_3_Left_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_3_Left_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_3_Left_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_3_Left_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_3_Left_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_3_Left_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_3_Left_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_3_Left_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_3_Left_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_3_Left_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_3_Left_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_3_Left_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_3_Left_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_3_Left_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_3_Left_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_3_Left_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_3_Left_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_3_Left_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_3_Left_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_3_Left_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_3_Left_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_3_Left_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_3_Left_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_3_Left_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_3_Left_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_3_Left_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_3_Left_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_3_Left_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_3_Left_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_3_Left_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_3_Left_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_3_Left_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_3_Left_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_3_Left_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_3_Left_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_3_Left_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_3_Left_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_3_Left_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_3_Left_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_3_Left_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_3_Left_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_3_Left_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_3_Left_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_3_Left_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_3_Left_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_3_Left_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_3_Left_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_3_Left_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_3_Left_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_3_Left_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_3_Left_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_3_Left_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_3_Left_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_3_Left_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_3_Left_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_3_Left_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_3_Left_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_3_Left_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_3_Left_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_3_Left_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_3_Left_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_3_Left_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_3_Left_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_3_Left_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_3_Left_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_3_Left_724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_3_Left_725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_3_Left_726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_3_Left_727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_3_Left_728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_3_Left_729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_3_Left_730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_3_Left_731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_3_Left_732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_3_Left_733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_3_Left_734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_3_Left_735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_3_Left_736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_3_Left_737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_3_Left_738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_3_Left_739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_3_Left_740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_3_Left_741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_3_Left_742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_3_Left_743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_3_Left_744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_3_Left_745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_3_Left_746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_3_Left_747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_3_Left_748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_3_Left_749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_3_Left_750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_3_Left_751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_3_Left_752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_3_Left_753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_3_Left_754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_3_Left_755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_3_Left_756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_3_Left_757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_3_Left_758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_3_Left_759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_3_Left_760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_3_Left_761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_3_Left_762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_3_Left_763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_3_Left_764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_3_Left_765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_3_Left_766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_3_Left_767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_3_Left_768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_3_Left_769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_3_Left_770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_3_Left_771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_3_Left_772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_3_Left_773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_3_Left_774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_3_Left_775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_3_Left_776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_3_Left_777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_3_Left_778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_3_Left_779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_3_Left_780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_3_Left_781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_3_Left_782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_3_Left_783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_3_Left_784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_3_Left_785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_3_Left_786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_3_Left_787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_3_Left_788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_3_Left_789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_3_Left_790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_3_Left_791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_3_Left_792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_3_Left_793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_3_Left_794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_3_Left_795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_3_Left_796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_3_Left_797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_3_Left_798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_3_Left_799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_3_Left_800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_3_Left_801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_3_Left_802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_3_Left_803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_3_Left_804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_3_Left_805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_3_Left_806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_3_Left_807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_3_Left_808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_3_Left_809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_3_Left_810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_3_Left_811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_3_Left_812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_3_Left_813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_3_Left_814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_3_Left_815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_3_Left_816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_3_Left_817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_3_Left_818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_3_Left_819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_3_Left_820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_3_Left_821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_3_Left_822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_3_Left_823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_3_Left_824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_3_Left_825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_3_Left_826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_3_Left_827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_3_Left_828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_3_Left_829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_3_Left_830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_3_Left_831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_3_Left_832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_3_Left_833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_3_Left_834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_3_Left_835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_3_Left_836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_3_Left_837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_3_Left_838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_3_Left_839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_3_Left_840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_3_Left_841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_3_Left_842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_3_Left_843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_3_Left_844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_3_Left_845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_3_Left_846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_3_Left_847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_3_Left_848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_3_Left_849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_3_Left_850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_3_Left_851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_3_Left_852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_3_Left_853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_3_Left_854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_3_Left_855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_3_Left_856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_3_Left_857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_3_Left_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_3_Left_859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_3_Left_860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_3_Left_861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_3_Left_862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_3_Left_863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_3_Left_864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_3_Left_865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_3_Left_866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_3_Left_867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_3_Left_868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_3_Left_869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_3_Left_870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_3_Left_871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_3_Left_872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_3_Left_873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_3_Left_874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_3_Left_875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_3_Left_876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_3_Left_877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_3_Left_878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_3_Left_879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_3_Left_880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_3_Left_881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_3_Left_882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_3_Left_883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_3_Left_884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_3_Left_885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_3_Left_886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_3_Left_887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_3_Left_888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_3_Left_889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_3_Left_890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_3_Left_891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_3_Left_892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_3_Left_893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_3_Left_894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_3_Left_895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_3_Left_896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_3_Left_897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_3_Left_898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_3_Left_899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_3_Left_900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_3_Left_901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_3_Left_902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_3_Left_903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_3_Left_904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_3_Left_905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_3_Left_906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_3_Left_907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_3_Left_908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_3_Left_909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_3_Left_910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_3_Left_911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_3_Left_912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_3_Left_913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_3_Left_914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_3_Left_915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_3_Left_916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_3_Left_917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_3_Left_918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_3_Left_919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_3_Left_920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_3_Left_921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_3_Left_922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_3_Left_923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_3_Left_924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_3_Left_925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_3_Left_926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_3_Left_927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_3_Left_928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_3_Left_929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_3_Left_930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_3_Left_931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_3_Left_932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_3_Left_933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_3_Left_934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_3_Left_935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_3_Left_936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_3_Left_937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_3_Left_938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_3_Left_939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_3_Left_940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_3_Left_941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_3_Left_942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_3_Left_943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_3_Left_944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_3_Left_945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_3_Left_946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_3_Left_947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_3_Left_948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_3_Left_949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_3_Left_950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_3_Left_951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_3_Left_952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_3_Left_953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_3_Left_954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_3_Left_955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_3_Left_956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_3_Left_957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_3_Left_958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_3_Left_959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_3_Left_960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_3_Left_961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_3_Left_962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_3_Left_963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_3_Left_964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_3_Left_965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_3_Left_966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_3_Left_967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_3_Left_968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_3_Left_969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_3_Left_970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_3_Left_971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_3_Right_972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_3_Right_973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_3_Right_974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_3_Right_975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_3_Right_976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_3_Right_977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_3_Right_978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_3_Right_979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_3_Right_980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_3_Right_981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_3_Right_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_3_Right_983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_3_Right_984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_3_Right_985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_3_Right_986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_3_Right_987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_3_Right_988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_3_Right_989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_3_Right_990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_3_Right_991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_3_Right_992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_3_Right_993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_3_Right_994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_3_Right_995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_3_Right_996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_3_Right_997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_3_Right_998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_3_Right_999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_3_Right_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_3_Right_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_3_Right_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_3_Right_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_3_Right_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_3_Right_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_3_Right_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_3_Right_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_3_Right_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_3_Right_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_3_Right_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_3_Right_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_3_Right_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_3_Right_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_3_Right_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_3_Right_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_3_Right_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_3_Right_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_3_Right_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_3_Right_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_3_Right_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_3_Right_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_3_Right_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_3_Right_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_3_Right_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_3_Right_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_3_Right_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_3_Right_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_3_Right_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_3_Right_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_3_Right_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_3_Right_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_3_Right_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_3_Right_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_3_Right_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_3_Right_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_3_Right_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_3_Right_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_3_Right_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_3_Right_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_3_Right_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_3_Right_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_3_Right_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_3_Right_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_3_Right_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_3_Right_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_3_Right_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_3_Right_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_3_Right_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_3_Right_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_3_Right_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_3_Right_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_3_Right_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_3_Right_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_3_Right_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_3_Right_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_3_Right_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_3_Right_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_3_Right_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_3_Right_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_3_Right_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_3_Right_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_3_Right_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_3_Right_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_3_Right_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_3_Right_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_3_Right_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_3_Right_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_3_Right_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_3_Right_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_3_Right_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_3_Right_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_3_Right_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_3_Right_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_3_Right_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_3_Right_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_3_Right_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_3_Right_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_3_Right_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_3_Right_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_3_Right_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_3_Right_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_3_Right_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_3_Right_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_3_Right_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_3_Right_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_3_Right_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_3_Right_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_3_Right_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_3_Right_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_3_Right_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_3_Right_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_3_Right_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_3_Right_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_3_Right_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_3_Right_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_3_Right_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_3_Right_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_3_Right_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_3_Right_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_3_Right_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_3_Right_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_3_Right_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_3_Right_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_3_Right_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_3_Right_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_3_Right_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_3_Right_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_3_Right_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_3_Right_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_3_Right_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_3_Right_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_3_Right_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_3_Right_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_3_Right_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_3_Right_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_3_Right_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_3_Right_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_3_Right_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_3_Right_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_3_Right_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_3_Right_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_3_Right_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_3_Right_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_3_Right_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_3_Right_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_3_Right_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_3_Right_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_3_Right_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_3_Right_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_3_Right_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_3_Right_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_3_Right_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_3_Right_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_3_Right_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_3_Right_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_3_Right_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_3_Right_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_3_Right_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_3_Right_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_3_Right_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_3_Right_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_3_Right_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_3_Right_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_3_Right_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_3_Right_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_3_Right_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_3_Right_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_3_Right_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_3_Right_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_3_Right_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_3_Right_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_3_Right_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_3_Right_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_3_Right_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_3_Right_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_3_Right_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_3_Right_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_3_Right_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_3_Right_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_3_Right_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_3_Right_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_3_Right_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_3_Right_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_3_Right_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_3_Right_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_3_Right_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_3_Right_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_3_Right_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_3_Right_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_3_Right_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_3_Right_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_3_Right_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_3_Right_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_3_Right_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_3_Right_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_3_Right_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_3_Right_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_3_Right_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_3_Right_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_3_Right_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_3_Right_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_3_Right_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_3_Right_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_3_Right_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_3_Right_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_3_Right_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_3_Right_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_3_Right_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_3_Right_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_3_Right_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_3_Right_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_3_Right_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_3_Right_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_3_Right_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_3_Right_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_3_Right_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_3_Right_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_3_Right_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_3_Right_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_3_Right_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_3_Right_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_3_Right_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_3_Right_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_3_Right_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_3_Right_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_3_Right_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_3_Right_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_3_Right_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_3_Right_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_3_Right_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_3_Right_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_3_Right_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_3_Right_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_3_Right_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_3_Right_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_3_Right_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_3_Right_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_3_Right_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_3_Right_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_3_Right_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_3_Right_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_3_Right_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_3_Right_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_3_Right_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_3_Right_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_3_Right_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_3_Right_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_3_Right_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_3_Right_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_3_Right_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_3_Right_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_3_Right_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_3_Right_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_3_Right_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_3_Right_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_3_Right_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_3_Right_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_3_Right_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_3_Right_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_3_Right_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_3_Right_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_3_Right_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_3_Right_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_3_Right_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_3_Right_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_3_Right_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_3_Right_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_3_Right_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_3_Right_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_3_Right_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_3_Right_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_3_Right_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_3_Right_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_3_Right_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_3_Right_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_3_Right_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_3_Right_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_3_Right_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_3_Right_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_3_Right_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_3_Right_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_3_Right_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_3_Right_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_3_Right_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_3_Right_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_3_Right_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_3_Right_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_3_Right_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_3_Right_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_3_Right_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_3_Right_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_3_Right_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_3_Right_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_3_Right_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_3_Right_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_3_Right_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_3_Right_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_3_Right_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_3_Right_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_3_Right_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_3_Right_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_3_Right_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_3_Right_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_3_Right_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_3_Right_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_3_Right_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_3_Right_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_3_Right_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_3_Right_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_3_Right_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_3_Right_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_3_Right_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_3_Right_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_3_Right_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_3_Right_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_4_Left_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_4_Left_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_4_Left_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_4_Left_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_4_Left_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_4_Left_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_4_Left_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_4_Left_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_4_Left_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_4_Left_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_4_Left_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_4_Left_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_4_Left_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_4_Left_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_4_Left_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_4_Left_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_4_Left_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_4_Left_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_4_Left_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_4_Left_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_4_Left_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_4_Left_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_4_Left_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_4_Left_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_4_Left_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_4_Left_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_4_Left_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_4_Left_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_4_Left_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_4_Left_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_4_Left_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_4_Left_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_4_Left_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_4_Left_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_4_Left_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_4_Left_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_4_Left_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_4_Left_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_4_Left_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_4_Left_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_4_Left_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_4_Left_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_4_Left_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_4_Left_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_4_Left_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_4_Left_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_4_Left_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_4_Left_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_4_Left_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_4_Left_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_4_Left_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_4_Left_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_4_Left_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_4_Left_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_4_Left_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_4_Left_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_4_Left_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_4_Left_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_4_Left_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_4_Left_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_4_Left_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_4_Left_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_4_Left_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_4_Left_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_4_Left_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_4_Left_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_4_Left_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_4_Left_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_4_Left_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_4_Left_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_4_Left_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_4_Left_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_4_Left_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_4_Left_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_4_Left_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_4_Left_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_4_Left_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_4_Left_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_4_Left_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_4_Left_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_4_Left_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_4_Left_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_4_Left_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_4_Left_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_4_Left_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_4_Left_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_4_Left_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_4_Left_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_4_Left_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_4_Left_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_4_Left_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_4_Left_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_4_Left_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_4_Left_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_4_Left_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_4_Left_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_4_Left_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_4_Left_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_4_Left_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_4_Left_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_4_Left_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_4_Left_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_4_Left_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_4_Left_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_4_Left_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_4_Left_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_4_Left_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_4_Left_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_4_Left_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_4_Left_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_4_Left_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_4_Left_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_4_Left_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_4_Left_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_4_Left_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_4_Left_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_4_Left_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_4_Left_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_4_Left_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_4_Left_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_4_Left_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_4_Left_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_4_Left_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_4_Left_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_4_Left_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_4_Left_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_4_Left_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_4_Left_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_4_Left_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_4_Left_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_4_Left_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_4_Left_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_4_Left_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_4_Left_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_4_Left_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_4_Left_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_4_Left_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_4_Left_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_4_Left_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_4_Left_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_4_Left_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_4_Left_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_4_Left_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_4_Left_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_4_Left_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_4_Left_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_4_Left_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_4_Left_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_4_Left_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_4_Left_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_4_Left_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_4_Left_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_4_Left_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_4_Left_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_4_Left_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_4_Left_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_4_Left_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_4_Left_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_4_Left_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_4_Left_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_4_Left_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_4_Left_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_4_Left_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_4_Left_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_4_Left_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_4_Left_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_4_Left_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_4_Left_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_4_Left_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_4_Left_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_4_Left_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_4_Left_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_4_Left_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_4_Left_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_4_Left_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_4_Left_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_4_Left_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_4_Left_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_4_Left_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_4_Left_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_4_Left_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_4_Left_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_4_Left_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_4_Left_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_4_Left_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_4_Left_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_4_Left_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_4_Left_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_4_Left_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_4_Left_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_4_Left_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_4_Left_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_4_Left_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_4_Left_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_4_Left_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_4_Left_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_4_Left_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_4_Left_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_4_Left_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_4_Left_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_4_Left_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_4_Left_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_4_Left_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_4_Left_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_4_Left_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_4_Left_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_4_Left_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_4_Left_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_4_Left_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_4_Left_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_4_Left_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_4_Left_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_4_Left_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_4_Left_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_4_Left_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_4_Left_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_4_Left_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_4_Left_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_4_Left_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_4_Left_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_4_Left_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_4_Left_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_4_Left_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_4_Left_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_4_Left_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_4_Left_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_4_Left_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_4_Left_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_4_Left_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_4_Left_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_4_Left_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_4_Left_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_4_Left_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_4_Left_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_4_Left_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_4_Left_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_4_Left_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_4_Left_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_4_Left_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_4_Left_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_4_Left_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_4_Left_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_4_Left_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_4_Left_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_4_Left_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_4_Left_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_4_Left_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_4_Left_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_4_Left_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_4_Left_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_4_Left_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_4_Left_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_4_Left_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_4_Left_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_4_Left_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_4_Left_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_4_Left_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_4_Left_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_4_Left_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_4_Left_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_4_Left_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_4_Left_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_4_Left_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_4_Left_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_4_Left_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_4_Left_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_4_Left_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_4_Left_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_4_Left_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_4_Left_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_4_Left_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_4_Left_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_4_Left_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_4_Left_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_4_Left_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_4_Left_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_4_Left_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_4_Left_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_4_Left_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_4_Left_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_4_Left_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_4_Left_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_4_Left_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_4_Left_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_4_Left_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_4_Left_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_4_Left_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_4_Left_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_4_Left_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_4_Left_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_4_Left_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_4_Left_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_4_Left_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_4_Left_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_4_Left_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_4_Left_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_4_Left_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_4_Left_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_4_Left_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_4_Left_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_4_Left_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_4_Left_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_4_Left_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_4_Left_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_4_Left_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_4_Left_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_4_Left_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_4_Left_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_4_Left_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_4_Left_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_4_Left_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_4_Left_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_4_Left_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_4_Left_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_4_Left_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_4_Left_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_4_Left_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_4_Left_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_4_Left_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_4_Left_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_4_Left_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_4_Left_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_4_Left_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_4_Left_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_4_Right_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_4_Right_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_4_Right_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_4_Right_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_4_Right_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_4_Right_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_4_Right_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_4_Right_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_4_Right_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_4_Right_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_4_Right_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_4_Right_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_4_Right_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_4_Right_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_4_Right_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_4_Right_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_4_Right_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_4_Right_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_4_Right_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_4_Right_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_4_Right_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_4_Right_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_4_Right_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_4_Right_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_4_Right_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_4_Right_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_4_Right_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_4_Right_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_4_Right_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_4_Right_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_4_Right_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_4_Right_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_4_Right_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_4_Right_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_4_Right_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_4_Right_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_4_Right_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_4_Right_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_4_Right_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_4_Right_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_4_Right_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_4_Right_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_4_Right_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_4_Right_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_4_Right_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_4_Right_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_4_Right_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_4_Right_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_4_Right_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_4_Right_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_4_Right_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_4_Right_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_4_Right_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_4_Right_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_4_Right_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_4_Right_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_4_Right_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_4_Right_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_4_Right_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_4_Right_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_4_Right_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_4_Right_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_4_Right_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_4_Right_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_4_Right_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_4_Right_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_4_Right_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_4_Right_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_4_Right_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_4_Right_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_4_Right_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_4_Right_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_4_Right_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_4_Right_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_4_Right_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_4_Right_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_4_Right_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_4_Right_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_4_Right_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_4_Right_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_4_Right_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_4_Right_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_4_Right_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_4_Right_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_4_Right_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_4_Right_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_4_Right_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_4_Right_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_4_Right_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_4_Right_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_4_Right_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_4_Right_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_4_Right_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_4_Right_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_4_Right_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_4_Right_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_4_Right_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_4_Right_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_4_Right_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_4_Right_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_4_Right_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_4_Right_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_4_Right_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_4_Right_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_4_Right_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_4_Right_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_4_Right_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_4_Right_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_4_Right_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_4_Right_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_4_Right_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_4_Right_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_4_Right_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_4_Right_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_4_Right_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_4_Right_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_4_Right_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_4_Right_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_4_Right_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_4_Right_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_4_Right_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_4_Right_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_4_Right_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_4_Right_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_4_Right_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_4_Right_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_4_Right_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_4_Right_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_4_Right_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_4_Right_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_4_Right_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_4_Right_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_4_Right_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_4_Right_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_4_Right_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_4_Right_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_4_Right_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_4_Right_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_4_Right_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_4_Right_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_4_Right_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_4_Right_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_4_Right_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_4_Right_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_4_Right_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_4_Right_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_4_Right_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_4_Right_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_4_Right_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_4_Right_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_4_Right_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_4_Right_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_4_Right_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_4_Right_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_4_Right_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_4_Right_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_4_Right_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_4_Right_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_4_Right_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_4_Right_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_4_Right_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_4_Right_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_4_Right_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_4_Right_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_4_Right_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_4_Right_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_4_Right_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_4_Right_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_4_Right_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_4_Right_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_4_Right_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_4_Right_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_4_Right_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_4_Right_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_4_Right_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_4_Right_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_4_Right_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_4_Right_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_4_Right_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_4_Right_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_4_Right_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_4_Right_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_4_Right_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_4_Right_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_4_Right_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_4_Right_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_4_Right_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_4_Right_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_4_Right_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_4_Right_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_4_Right_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_4_Right_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_4_Right_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_4_Right_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_4_Right_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_4_Right_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_4_Right_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_4_Right_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_4_Right_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_4_Right_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_4_Right_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_4_Right_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_4_Right_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_4_Right_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_4_Right_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_4_Right_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_4_Right_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_4_Right_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_4_Right_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_4_Right_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_4_Right_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_4_Right_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_4_Right_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_4_Right_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_4_Right_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_4_Right_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_4_Right_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_4_Right_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_4_Right_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_4_Right_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_4_Right_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_4_Right_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_4_Right_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_4_Right_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_4_Right_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_4_Right_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_4_Right_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_4_Right_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_4_Right_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_4_Right_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_4_Right_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_4_Right_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_4_Right_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_4_Right_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_4_Right_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_4_Right_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_4_Right_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_4_Right_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_4_Right_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_4_Right_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_4_Right_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_4_Right_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_4_Right_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_4_Right_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_4_Right_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_4_Right_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_4_Right_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_4_Right_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_4_Right_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_4_Right_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_4_Right_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_4_Right_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_4_Right_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_4_Right_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_4_Right_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_4_Right_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_4_Right_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_4_Right_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_4_Right_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_4_Right_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_4_Right_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_4_Right_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_4_Right_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_4_Right_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_4_Right_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_4_Right_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_4_Right_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_4_Right_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_4_Right_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_4_Right_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_4_Right_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_4_Right_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_4_Right_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_4_Right_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_4_Right_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_4_Right_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_4_Right_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_4_Right_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_4_Right_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_4_Right_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_4_Right_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_4_Right_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_4_Right_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_4_Right_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_4_Right_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_4_Right_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_4_Right_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_4_Right_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_4_Right_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_4_Right_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_4_Right_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_4_Right_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_4_Right_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_4_Right_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_4_Right_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_4_Right_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_4_Right_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_4_Right_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_4_Right_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_4_Right_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_4_Right_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_4_Right_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_4_Right_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_4_Right_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_4_Right_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_4_Right_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_4_Right_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_4_Right_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_4_Right_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_4_Right_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_4_Right_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_4_Right_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_4_Right_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_4_Right_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_4_Right_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_4_Right_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_4_Right_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_4_Right_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_4_Right_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_4_Right_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_4_Right_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_4_Right_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_4_Right_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_4_Right_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_5_Left_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_5_Left_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_5_Left_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_5_Left_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_5_Left_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_5_Left_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_5_Left_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_5_Left_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_5_Left_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_5_Left_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_5_Left_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_5_Left_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_5_Left_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_5_Left_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_5_Left_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_5_Left_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_5_Left_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_5_Left_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_5_Left_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_5_Left_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_5_Left_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_5_Left_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_5_Left_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_5_Left_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_5_Left_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_5_Left_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_5_Left_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_5_Left_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_5_Left_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_5_Left_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_5_Left_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_5_Left_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_5_Left_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_5_Left_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_5_Left_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_5_Left_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_5_Left_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_5_Left_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_5_Left_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_5_Left_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_5_Left_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_5_Left_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_5_Left_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_5_Left_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_5_Left_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_5_Left_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_5_Left_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_5_Left_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_5_Left_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_5_Left_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_5_Left_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_5_Left_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_5_Left_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_5_Left_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_5_Left_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_5_Left_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_5_Left_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_5_Left_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_5_Left_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_5_Left_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_5_Left_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_5_Left_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_5_Left_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_5_Left_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_5_Left_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_5_Left_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_5_Left_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_5_Left_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_5_Left_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_5_Left_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_5_Left_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_5_Left_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_5_Left_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_5_Left_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_5_Left_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_5_Left_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_5_Left_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_5_Left_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_5_Left_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_5_Left_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_5_Left_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_5_Left_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_5_Left_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_5_Left_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_5_Left_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_5_Left_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_5_Left_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_5_Left_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_5_Left_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_5_Left_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_5_Left_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_5_Left_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_5_Left_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_5_Left_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_5_Left_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_5_Left_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_5_Left_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_5_Left_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_5_Left_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_5_Left_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_5_Left_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_5_Left_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_5_Left_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_5_Left_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_5_Left_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_5_Left_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_5_Left_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_5_Left_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_5_Left_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_5_Left_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_5_Left_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_5_Left_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_5_Left_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_5_Left_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_5_Left_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_5_Left_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_5_Left_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_5_Left_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_5_Left_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_5_Left_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_5_Left_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_5_Left_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_5_Left_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_5_Left_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_5_Left_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_5_Left_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_5_Left_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_5_Left_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_5_Left_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_5_Left_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_5_Left_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_5_Left_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_5_Left_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_5_Left_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_5_Left_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_5_Left_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_5_Left_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_5_Left_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_5_Left_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_5_Left_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_5_Left_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_5_Left_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_5_Left_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_5_Left_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_5_Left_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_5_Left_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_5_Left_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_5_Left_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_5_Left_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_5_Left_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_5_Left_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_5_Left_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_5_Left_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_5_Left_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_5_Left_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_5_Left_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_5_Left_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_5_Left_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_5_Left_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_5_Left_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_5_Left_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_5_Left_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_5_Left_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_5_Left_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_5_Left_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_5_Left_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_5_Left_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_5_Left_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_5_Left_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_5_Left_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_5_Left_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_5_Left_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_5_Left_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_5_Left_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_5_Left_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_5_Left_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_5_Left_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_5_Left_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_5_Left_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_5_Left_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_5_Left_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_5_Left_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_5_Left_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_5_Left_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_5_Left_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_5_Left_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_5_Left_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_5_Left_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_5_Left_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_5_Left_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_5_Left_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_5_Left_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_5_Left_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_5_Left_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_5_Left_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_5_Left_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_5_Left_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_5_Left_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_5_Left_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_5_Left_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_5_Left_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_5_Left_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_5_Left_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_5_Left_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_5_Left_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_5_Left_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_5_Left_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_5_Left_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_5_Left_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_5_Left_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_5_Left_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_5_Left_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_5_Left_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_5_Left_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_5_Left_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_5_Left_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_5_Left_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_5_Left_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_5_Left_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_5_Left_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_5_Left_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_5_Left_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_5_Left_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_5_Left_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_5_Left_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_5_Left_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_5_Left_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_5_Left_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_5_Left_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_5_Left_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_5_Left_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_5_Left_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_5_Left_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_5_Left_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_5_Left_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_5_Left_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_5_Left_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_5_Left_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_5_Left_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_5_Left_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_5_Left_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_5_Left_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_5_Left_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_5_Left_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_5_Left_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_5_Left_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_5_Left_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_5_Left_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_5_Left_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_5_Left_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_5_Left_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_5_Left_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_5_Left_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_5_Left_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_5_Left_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_5_Left_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_5_Left_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_5_Left_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_5_Left_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_5_Left_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_5_Left_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_5_Left_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_5_Left_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_5_Left_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_5_Left_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_5_Left_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_5_Left_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_5_Left_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_5_Left_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_5_Left_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_5_Left_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_5_Left_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_5_Left_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_5_Left_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_5_Left_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_5_Left_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_5_Left_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_5_Left_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_5_Left_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_5_Left_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_5_Left_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_5_Left_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_5_Left_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_5_Left_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_5_Left_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_5_Left_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_5_Left_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_5_Left_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_5_Left_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_5_Left_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_5_Left_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_5_Left_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_5_Left_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_5_Left_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_5_Left_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_5_Left_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_5_Left_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_5_Left_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_5_Left_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_5_Left_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_5_Left_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_5_Left_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_5_Left_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_5_Left_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_5_Left_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_5_Left_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_5_Left_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_5_Left_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_5_Left_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_5_Left_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_5_Left_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_5_Left_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_5_Left_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_5_Left_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_5_Left_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_5_Left_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_5_Left_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_5_Left_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_5_Left_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_5_Left_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_5_Left_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_5_Left_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_5_Left_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_5_Left_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_5_Right_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_5_Right_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_5_Right_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_5_Right_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_5_Right_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_5_Right_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_5_Right_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_5_Right_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_5_Right_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_5_Right_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_5_Right_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_5_Right_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_5_Right_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_5_Right_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_5_Right_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_5_Right_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_5_Right_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_5_Right_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_5_Right_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_5_Right_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_5_Right_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_5_Right_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_5_Right_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_5_Right_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_5_Right_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_5_Right_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_5_Right_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_5_Right_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_5_Right_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_5_Right_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_5_Right_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_5_Right_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_5_Right_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_5_Right_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_5_Right_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_5_Right_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_5_Right_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_5_Right_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_5_Right_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_5_Right_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_5_Right_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_5_Right_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_5_Right_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_5_Right_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_5_Right_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_5_Right_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_5_Right_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_5_Right_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_5_Right_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_5_Right_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_5_Right_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_5_Right_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_5_Right_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_5_Right_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_5_Right_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_5_Right_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_5_Right_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_5_Right_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_5_Right_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_5_Right_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_5_Right_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_5_Right_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_5_Right_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_5_Right_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_5_Right_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_5_Right_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_5_Right_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_5_Right_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_5_Right_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_5_Right_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_5_Right_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_5_Right_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_5_Right_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_5_Right_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_5_Right_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_5_Right_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_5_Right_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_5_Right_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_5_Right_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_5_Right_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_5_Right_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_5_Right_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_5_Right_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_5_Right_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_5_Right_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_5_Right_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_5_Right_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_5_Right_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_5_Right_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_5_Right_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_5_Right_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_5_Right_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_5_Right_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_5_Right_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_5_Right_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_5_Right_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_5_Right_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_5_Right_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_5_Right_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_5_Right_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_5_Right_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_5_Right_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_5_Right_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_5_Right_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_5_Right_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_5_Right_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_5_Right_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_5_Right_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_5_Right_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_5_Right_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_5_Right_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_5_Right_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_5_Right_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_5_Right_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_5_Right_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_5_Right_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_5_Right_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_5_Right_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_5_Right_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_5_Right_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_5_Right_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_5_Right_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_5_Right_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_5_Right_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_5_Right_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_5_Right_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_5_Right_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_5_Right_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_5_Right_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_5_Right_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_5_Right_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_5_Right_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_5_Right_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_5_Right_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_5_Right_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_5_Right_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_5_Right_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_5_Right_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_5_Right_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_5_Right_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_5_Right_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_5_Right_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_5_Right_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_5_Right_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_5_Right_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_5_Right_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_5_Right_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_5_Right_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_5_Right_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_5_Right_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_5_Right_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_5_Right_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_5_Right_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_5_Right_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_5_Right_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_5_Right_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_5_Right_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_5_Right_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_5_Right_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_5_Right_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_5_Right_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_5_Right_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_5_Right_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_5_Right_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_5_Right_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_5_Right_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_5_Right_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_5_Right_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_5_Right_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_5_Right_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_5_Right_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_5_Right_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_5_Right_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_5_Right_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_5_Right_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_5_Right_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_5_Right_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_5_Right_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_5_Right_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_5_Right_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_5_Right_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_5_Right_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_5_Right_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_5_Right_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_5_Right_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_5_Right_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_5_Right_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_5_Right_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_5_Right_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_5_Right_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_5_Right_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_5_Right_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_5_Right_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_5_Right_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_5_Right_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_5_Right_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_5_Right_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_5_Right_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_5_Right_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_5_Right_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_5_Right_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_5_Right_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_5_Right_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_5_Right_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_5_Right_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_5_Right_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_5_Right_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_5_Right_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_5_Right_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_5_Right_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_5_Right_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_5_Right_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_5_Right_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_5_Right_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_5_Right_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_5_Right_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_5_Right_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_5_Right_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_5_Right_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_5_Right_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_5_Right_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_5_Right_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_5_Right_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_5_Right_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_5_Right_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_5_Right_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_5_Right_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_5_Right_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_5_Right_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_5_Right_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_5_Right_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_5_Right_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_5_Right_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_5_Right_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_5_Right_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_5_Right_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_5_Right_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_5_Right_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_5_Right_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_5_Right_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_5_Right_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_5_Right_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_5_Right_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_5_Right_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_5_Right_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_5_Right_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_5_Right_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_5_Right_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_5_Right_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_5_Right_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_5_Right_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_5_Right_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_5_Right_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_5_Right_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_5_Right_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_5_Right_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_5_Right_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_5_Right_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_5_Right_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_5_Right_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_5_Right_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_5_Right_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_5_Right_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_5_Right_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_5_Right_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_5_Right_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_5_Right_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_5_Right_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_5_Right_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_5_Right_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_5_Right_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_5_Right_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_5_Right_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_5_Right_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_5_Right_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_5_Right_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_5_Right_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_5_Right_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_5_Right_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_5_Right_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_5_Right_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_5_Right_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_5_Right_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_5_Right_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_5_Right_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_5_Right_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_5_Right_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_5_Right_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_5_Right_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_5_Right_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_5_Right_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_5_Right_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_5_Right_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_5_Right_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_5_Right_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_5_Right_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_5_Right_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_5_Right_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_5_Right_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_5_Right_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_5_Right_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_5_Right_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_5_Right_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_5_Right_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_5_Right_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_5_Right_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_5_Right_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_5_Right_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_5_Right_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_5_Right_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_5_Right_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_5_Right_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_5_Right_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_5_Right_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_5_Right_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_5_Right_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_5_Right_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_5_Right_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_5_Right_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_5_Right_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_5_Right_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_5_Right_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_5_Right_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_5_Right_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_6_Left_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_6_Left_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_6_Left_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_6_Left_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_6_Left_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_6_Left_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_6_Left_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_6_Left_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_6_Left_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_6_Left_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_6_Left_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_6_Left_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_6_Left_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_6_Left_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_6_Left_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_6_Left_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_6_Left_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_6_Left_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_6_Left_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_6_Left_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_6_Left_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_6_Left_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_6_Left_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_6_Left_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_6_Left_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_6_Left_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_6_Left_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_6_Left_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_6_Left_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_6_Left_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_6_Left_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_6_Left_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_6_Left_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_6_Left_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_6_Left_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_6_Left_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_6_Left_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_6_Left_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_6_Left_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_6_Left_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_6_Left_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_6_Left_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_6_Left_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_6_Left_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_6_Left_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_6_Left_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_6_Left_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_6_Left_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_6_Left_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_6_Left_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_6_Left_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_6_Left_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_6_Left_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_6_Left_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_6_Left_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_6_Left_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_6_Left_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_6_Left_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_6_Left_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_6_Left_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_6_Left_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_6_Left_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_6_Left_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_6_Left_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_6_Left_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_6_Left_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_6_Left_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_6_Left_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_6_Left_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_6_Left_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_6_Left_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_6_Left_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_6_Left_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_6_Left_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_6_Left_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_6_Left_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_6_Left_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_6_Left_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_6_Left_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_6_Left_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_6_Left_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_6_Left_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_6_Left_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_6_Left_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_6_Left_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_6_Left_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_6_Left_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_6_Left_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_6_Left_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_6_Left_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_6_Left_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_6_Left_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_6_Left_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_6_Left_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_6_Left_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_6_Left_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_6_Left_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_6_Left_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_6_Left_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_6_Left_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_6_Left_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_6_Left_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_6_Left_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_6_Left_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_6_Left_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_6_Left_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_6_Left_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_6_Left_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_6_Left_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_6_Left_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_6_Left_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_6_Left_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_6_Left_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_6_Left_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_6_Left_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_6_Left_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_6_Left_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_6_Left_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_6_Left_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_6_Left_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_6_Left_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_6_Left_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_6_Left_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_6_Left_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_6_Left_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_6_Left_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_6_Left_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_6_Left_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_6_Left_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_6_Left_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_6_Left_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_6_Left_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_6_Left_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_6_Left_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_6_Left_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_6_Left_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_6_Left_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_6_Left_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_6_Left_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_6_Left_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_6_Left_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_6_Left_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_6_Left_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_6_Left_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_6_Left_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_6_Left_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_6_Left_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_6_Left_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_6_Left_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_6_Left_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_6_Left_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_6_Left_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_6_Left_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_6_Left_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_6_Left_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_6_Left_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_6_Left_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_6_Left_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_6_Left_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_6_Left_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_6_Left_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_6_Left_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_6_Left_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_6_Left_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_6_Left_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_6_Left_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_6_Left_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_6_Left_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_6_Left_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_6_Left_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_6_Left_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_6_Left_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_6_Left_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_6_Left_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_6_Left_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_6_Left_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_6_Left_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_6_Left_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_6_Left_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_6_Left_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_6_Left_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_6_Left_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_6_Left_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_6_Left_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_6_Left_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_6_Left_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_6_Left_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_6_Left_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_6_Left_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_6_Left_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_6_Left_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_6_Left_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_6_Left_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_6_Left_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_6_Left_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_6_Left_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_6_Left_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_6_Left_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_6_Left_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_6_Left_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_6_Left_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_6_Left_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_6_Left_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_6_Left_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_6_Left_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_6_Left_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_6_Left_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_6_Left_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_6_Left_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_6_Left_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_6_Left_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_6_Left_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_6_Left_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_6_Left_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_6_Left_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_6_Left_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_6_Left_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_6_Left_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_6_Left_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_6_Left_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_6_Left_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_6_Left_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_6_Left_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_6_Left_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_6_Left_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_6_Left_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_6_Left_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_6_Left_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_6_Left_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_6_Left_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_6_Left_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_6_Left_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_6_Left_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_6_Left_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_6_Left_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_6_Left_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_6_Left_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_6_Left_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_6_Left_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_6_Left_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_6_Left_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_6_Left_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_6_Left_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_6_Left_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_6_Left_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_6_Left_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_6_Left_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_6_Left_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_6_Left_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_6_Left_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_6_Left_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_6_Left_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_6_Left_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_6_Left_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_6_Left_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_6_Left_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_6_Left_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_6_Left_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_6_Left_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_6_Left_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_6_Left_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_6_Left_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_6_Left_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_6_Left_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_6_Left_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_6_Left_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_6_Left_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_6_Left_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_6_Left_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_6_Left_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_6_Left_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_6_Left_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_6_Left_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_6_Left_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_6_Left_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_6_Left_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_6_Left_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_6_Left_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_6_Left_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_6_Left_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_6_Left_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_6_Left_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_6_Left_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_6_Left_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_6_Left_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_6_Left_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_6_Left_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_6_Left_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_6_Left_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_6_Left_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_6_Left_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_6_Left_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_6_Left_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_6_Left_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_6_Left_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_6_Left_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_6_Left_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_6_Left_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_6_Left_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_6_Left_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_6_Left_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_6_Left_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_6_Left_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_6_Left_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_6_Left_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_6_Left_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_6_Left_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_6_Left_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_6_Left_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_6_Left_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_6_Left_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_6_Left_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_6_Left_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_6_Left_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_6_Left_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_6_Left_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_6_Left_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_6_Left_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_6_Left_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_6_Left_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_6_Left_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_6_Left_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_6_Left_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_6_Left_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_6_Right_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_6_Right_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_6_Right_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_6_Right_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_6_Right_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_6_Right_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_6_Right_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_6_Right_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_6_Right_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_6_Right_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_6_Right_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_6_Right_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_6_Right_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_6_Right_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_6_Right_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_6_Right_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_6_Right_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_6_Right_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_6_Right_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_6_Right_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_6_Right_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_6_Right_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_6_Right_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_6_Right_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_6_Right_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_6_Right_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_6_Right_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_6_Right_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_6_Right_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_6_Right_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_6_Right_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_6_Right_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_6_Right_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_6_Right_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_6_Right_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_6_Right_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_6_Right_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_6_Right_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_6_Right_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_6_Right_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_6_Right_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_6_Right_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_6_Right_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_6_Right_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_6_Right_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_6_Right_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_6_Right_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_6_Right_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_6_Right_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_6_Right_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_6_Right_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_6_Right_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_6_Right_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_6_Right_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_6_Right_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_6_Right_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_6_Right_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_6_Right_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_6_Right_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_6_Right_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_6_Right_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_6_Right_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_6_Right_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_6_Right_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_6_Right_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_6_Right_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_6_Right_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_6_Right_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_6_Right_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_6_Right_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_6_Right_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_6_Right_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_6_Right_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_6_Right_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_6_Right_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_6_Right_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_6_Right_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_6_Right_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_6_Right_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_6_Right_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_6_Right_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_6_Right_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_6_Right_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_6_Right_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_6_Right_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_6_Right_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_6_Right_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_6_Right_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_6_Right_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_6_Right_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_6_Right_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_6_Right_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_6_Right_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_6_Right_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_6_Right_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_6_Right_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_6_Right_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_6_Right_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_6_Right_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_6_Right_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_6_Right_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_6_Right_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_6_Right_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_6_Right_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_6_Right_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_6_Right_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_6_Right_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_6_Right_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_6_Right_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_6_Right_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_6_Right_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_6_Right_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_6_Right_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_6_Right_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_6_Right_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_6_Right_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_6_Right_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_6_Right_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_6_Right_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_6_Right_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_6_Right_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_6_Right_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_6_Right_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_6_Right_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_6_Right_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_6_Right_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_6_Right_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_6_Right_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_6_Right_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_6_Right_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_6_Right_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_6_Right_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_6_Right_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_6_Right_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_6_Right_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_6_Right_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_6_Right_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_6_Right_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_6_Right_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_6_Right_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_6_Right_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_6_Right_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_6_Right_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_6_Right_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_6_Right_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_6_Right_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_6_Right_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_6_Right_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_6_Right_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_6_Right_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_6_Right_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_6_Right_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_6_Right_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_6_Right_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_6_Right_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_6_Right_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_6_Right_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_6_Right_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_6_Right_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_6_Right_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_6_Right_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_6_Right_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_6_Right_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_6_Right_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_6_Right_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_6_Right_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_6_Right_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_6_Right_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_6_Right_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_6_Right_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_6_Right_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_6_Right_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_6_Right_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_6_Right_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_6_Right_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_6_Right_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_6_Right_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_6_Right_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_6_Right_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_6_Right_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_6_Right_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_6_Right_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_6_Right_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_6_Right_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_6_Right_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_6_Right_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_6_Right_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_6_Right_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_6_Right_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_6_Right_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_6_Right_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_6_Right_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_6_Right_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_6_Right_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_6_Right_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_6_Right_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_6_Right_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_6_Right_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_6_Right_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_6_Right_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_6_Right_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_6_Right_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_6_Right_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_6_Right_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_6_Right_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_6_Right_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_6_Right_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_6_Right_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_6_Right_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_6_Right_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_6_Right_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_6_Right_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_6_Right_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_6_Right_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_6_Right_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_6_Right_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_6_Right_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_6_Right_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_6_Right_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_6_Right_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_6_Right_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_6_Right_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_6_Right_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_6_Right_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_6_Right_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_6_Right_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_6_Right_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_6_Right_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_6_Right_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_6_Right_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_6_Right_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_6_Right_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_6_Right_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_6_Right_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_6_Right_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_6_Right_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_6_Right_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_6_Right_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_6_Right_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_6_Right_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_6_Right_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_6_Right_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_6_Right_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_6_Right_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_6_Right_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_6_Right_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_6_Right_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_6_Right_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_6_Right_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_6_Right_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_6_Right_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_6_Right_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_6_Right_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_6_Right_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_6_Right_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_6_Right_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_6_Right_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_6_Right_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_6_Right_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_6_Right_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_6_Right_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_6_Right_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_6_Right_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_6_Right_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_6_Right_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_6_Right_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_6_Right_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_6_Right_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_6_Right_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_6_Right_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_6_Right_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_6_Right_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_6_Right_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_6_Right_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_6_Right_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_6_Right_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_6_Right_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_6_Right_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_6_Right_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_6_Right_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_6_Right_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_6_Right_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_6_Right_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_6_Right_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_6_Right_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_6_Right_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_6_Right_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_6_Right_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_6_Right_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_6_Right_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_6_Right_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_6_Right_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_6_Right_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_6_Right_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_6_Right_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_6_Right_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_6_Right_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_6_Right_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_6_Right_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_6_Right_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_6_Right_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_6_Right_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_6_Right_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_6_Right_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_6_Right_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_6_Right_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_6_Right_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_6_Right_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_6_Right_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_6_Right_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_6_Right_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_6_Right_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_6_Right_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_6_Right_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_6_Right_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_6_Right_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_6_Right_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_6_Right_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_6_Right_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_6_Right_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_6_Right_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_6_Right_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_6_Right_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_6_Right_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_7_Left_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_7_Left_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_7_Left_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_7_Left_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_7_Left_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_7_Left_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_7_Left_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_7_Left_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_7_Left_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_7_Left_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_7_Left_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_7_Left_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_7_Left_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_7_Left_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_7_Left_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_7_Left_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_7_Left_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_7_Left_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_7_Left_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_7_Left_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_7_Left_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_7_Left_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_7_Left_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_7_Left_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_7_Left_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_7_Left_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_7_Left_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_7_Left_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_7_Left_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_7_Left_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_7_Left_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_7_Left_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_7_Left_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_7_Left_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_7_Left_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_7_Left_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_7_Left_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_7_Left_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_7_Left_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_7_Left_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_7_Left_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_7_Left_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_7_Left_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_7_Left_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_7_Left_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_7_Left_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_7_Left_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_7_Left_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_7_Left_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_7_Left_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_7_Left_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_7_Left_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_7_Left_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_7_Left_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_7_Left_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_7_Left_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_7_Left_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_7_Left_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_7_Left_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_7_Left_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_7_Left_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_7_Left_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_7_Left_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_7_Left_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_7_Left_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_7_Left_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_7_Left_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_7_Left_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_7_Left_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_7_Left_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_7_Left_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_7_Left_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_7_Left_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_7_Left_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_7_Left_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_7_Left_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_7_Left_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_7_Left_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_7_Left_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_7_Left_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_7_Left_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_7_Left_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_7_Left_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_7_Left_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_7_Left_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_7_Left_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_7_Left_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_7_Left_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_7_Left_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_7_Left_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_7_Left_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_7_Left_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_7_Left_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_7_Left_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_7_Left_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_7_Left_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_7_Left_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_7_Left_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_7_Left_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_7_Left_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_7_Left_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_7_Left_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_7_Left_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_7_Left_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_7_Left_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_7_Left_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_7_Left_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_7_Left_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_7_Left_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_7_Left_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_7_Left_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_7_Left_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_7_Left_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_7_Left_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_7_Left_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_7_Left_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_7_Left_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_7_Left_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_7_Left_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_7_Left_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_7_Left_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_7_Left_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_7_Left_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_7_Left_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_7_Left_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_7_Left_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_7_Left_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_7_Left_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_7_Left_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_7_Left_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_7_Left_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_7_Left_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_7_Left_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_7_Left_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_7_Left_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_7_Left_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_7_Left_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_7_Left_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_7_Left_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_7_Left_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_7_Left_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_7_Left_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_7_Left_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_7_Left_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_7_Left_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_7_Left_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_7_Left_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_7_Left_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_7_Left_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_7_Left_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_7_Left_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_7_Left_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_7_Left_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_7_Left_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_7_Left_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_7_Left_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_7_Left_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_7_Left_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_7_Left_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_7_Left_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_7_Left_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_7_Left_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_7_Left_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_7_Left_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_7_Left_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_7_Left_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_7_Left_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_7_Left_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_7_Left_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_7_Left_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_7_Left_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_7_Left_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_7_Left_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_7_Left_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_7_Left_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_7_Left_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_7_Left_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_7_Left_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_7_Left_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_7_Left_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_7_Left_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_7_Left_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_7_Left_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_7_Left_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_7_Left_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_7_Left_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_7_Left_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_7_Left_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_7_Left_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_7_Left_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_7_Left_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_7_Left_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_7_Left_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_7_Left_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_7_Left_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_7_Left_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_7_Left_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_7_Left_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_7_Left_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_7_Left_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_7_Left_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_7_Left_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_7_Left_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_7_Left_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_7_Left_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_7_Left_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_7_Left_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_7_Left_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_7_Left_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_7_Left_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_7_Left_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_7_Left_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_7_Left_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_7_Left_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_7_Left_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_7_Left_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_7_Left_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_7_Left_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_7_Left_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_7_Left_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_7_Left_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_7_Left_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_7_Left_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_7_Left_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_7_Left_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_7_Left_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_7_Left_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_7_Left_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_7_Left_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_7_Left_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_7_Left_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_7_Left_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_7_Left_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_7_Left_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_7_Left_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_7_Left_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_7_Left_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_7_Left_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_7_Left_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_7_Left_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_7_Left_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_7_Left_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_7_Left_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_7_Left_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_7_Left_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_7_Left_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_7_Left_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_7_Left_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_7_Left_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_7_Left_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_7_Left_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_7_Left_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_7_Left_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_7_Left_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_7_Left_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_7_Left_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_7_Left_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_7_Left_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_7_Left_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_7_Left_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_7_Left_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_7_Left_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_7_Left_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_7_Left_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_7_Left_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_7_Left_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_7_Left_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_7_Left_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_7_Left_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_7_Left_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_7_Left_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_7_Left_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_7_Left_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_7_Left_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_7_Left_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_7_Left_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_7_Left_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_7_Left_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_7_Left_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_7_Left_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_7_Left_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_7_Left_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_7_Left_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_7_Left_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_7_Left_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_7_Left_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_7_Left_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_7_Left_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_7_Left_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_7_Left_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_7_Left_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_7_Left_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_7_Left_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_7_Left_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_7_Left_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_7_Left_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_7_Left_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_7_Left_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_7_Left_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_7_Left_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_7_Left_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_7_Left_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_7_Left_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_7_Left_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_7_Left_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_7_Left_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_7_Left_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_7_Left_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_7_Left_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_7_Left_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_7_Left_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_7_Left_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_7_Left_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_7_Left_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_7_Left_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_7_Left_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_7_Left_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_7_Left_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_7_Left_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_7_Left_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_7_Left_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_7_Left_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_7_Left_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_7_Left_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_7_Right_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_7_Right_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_7_Right_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_7_Right_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_7_Right_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_7_Right_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_7_Right_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_7_Right_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_7_Right_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_7_Right_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_7_Right_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_7_Right_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_7_Right_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_7_Right_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_7_Right_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_7_Right_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_7_Right_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_7_Right_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_7_Right_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_7_Right_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_7_Right_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_7_Right_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_7_Right_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_7_Right_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_7_Right_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_7_Right_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_7_Right_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_7_Right_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_7_Right_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_7_Right_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_7_Right_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_7_Right_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_7_Right_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_7_Right_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_7_Right_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_7_Right_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_7_Right_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_7_Right_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_7_Right_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_7_Right_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_7_Right_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_7_Right_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_7_Right_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_7_Right_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_7_Right_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_7_Right_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_7_Right_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_7_Right_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_7_Right_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_7_Right_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_7_Right_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_7_Right_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_7_Right_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_7_Right_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_7_Right_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_7_Right_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_7_Right_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_7_Right_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_7_Right_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_7_Right_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_7_Right_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_7_Right_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_7_Right_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_7_Right_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_7_Right_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_7_Right_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_7_Right_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_7_Right_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_7_Right_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_7_Right_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_7_Right_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_7_Right_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_7_Right_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_7_Right_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_7_Right_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_7_Right_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_7_Right_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_7_Right_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_7_Right_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_7_Right_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_7_Right_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_7_Right_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_7_Right_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_7_Right_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_7_Right_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_7_Right_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_7_Right_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_7_Right_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_7_Right_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_7_Right_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_7_Right_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_7_Right_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_7_Right_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_7_Right_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_7_Right_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_7_Right_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_7_Right_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_7_Right_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_7_Right_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_7_Right_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_7_Right_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_7_Right_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_7_Right_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_7_Right_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_7_Right_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_7_Right_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_7_Right_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_7_Right_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_7_Right_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_7_Right_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_7_Right_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_7_Right_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_7_Right_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_7_Right_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_7_Right_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_7_Right_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_7_Right_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_7_Right_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_7_Right_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_7_Right_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_7_Right_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_7_Right_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_7_Right_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_7_Right_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_7_Right_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_7_Right_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_7_Right_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_7_Right_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_7_Right_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_7_Right_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_7_Right_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_7_Right_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_7_Right_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_7_Right_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_7_Right_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_7_Right_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_7_Right_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_7_Right_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_7_Right_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_7_Right_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_7_Right_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_7_Right_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_7_Right_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_7_Right_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_7_Right_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_7_Right_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_7_Right_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_7_Right_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_7_Right_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_7_Right_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_7_Right_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_7_Right_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_7_Right_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_7_Right_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_7_Right_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_7_Right_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_7_Right_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_7_Right_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_7_Right_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_7_Right_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_7_Right_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_7_Right_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_7_Right_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_7_Right_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_7_Right_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_7_Right_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_7_Right_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_7_Right_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_7_Right_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_7_Right_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_7_Right_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_7_Right_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_7_Right_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_7_Right_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_7_Right_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_7_Right_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_7_Right_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_7_Right_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_7_Right_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_7_Right_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_7_Right_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_7_Right_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_7_Right_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_7_Right_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_7_Right_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_7_Right_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_7_Right_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_7_Right_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_7_Right_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_7_Right_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_7_Right_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_7_Right_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_7_Right_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_7_Right_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_7_Right_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_7_Right_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_7_Right_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_7_Right_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_7_Right_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_7_Right_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_7_Right_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_7_Right_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_7_Right_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_7_Right_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_7_Right_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_7_Right_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_7_Right_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_7_Right_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_7_Right_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_7_Right_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_7_Right_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_7_Right_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_7_Right_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_7_Right_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_7_Right_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_7_Right_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_7_Right_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_7_Right_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_7_Right_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_7_Right_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_7_Right_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_7_Right_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_7_Right_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_7_Right_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_7_Right_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_7_Right_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_7_Right_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_7_Right_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_7_Right_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_7_Right_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_7_Right_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_7_Right_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_7_Right_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_7_Right_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_7_Right_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_7_Right_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_7_Right_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_7_Right_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_7_Right_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_7_Right_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_7_Right_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_7_Right_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_7_Right_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_7_Right_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_7_Right_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_7_Right_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_7_Right_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_7_Right_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_7_Right_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_7_Right_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_7_Right_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_7_Right_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_7_Right_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_7_Right_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_7_Right_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_7_Right_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_7_Right_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_7_Right_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_7_Right_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_7_Right_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_7_Right_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_7_Right_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_7_Right_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_7_Right_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_7_Right_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_7_Right_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_7_Right_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_7_Right_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_7_Right_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_7_Right_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_7_Right_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_7_Right_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_7_Right_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_7_Right_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_7_Right_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_7_Right_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_7_Right_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_7_Right_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_7_Right_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_7_Right_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_7_Right_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_7_Right_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_7_Right_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_7_Right_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_7_Right_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_7_Right_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_7_Right_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_7_Right_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_7_Right_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_7_Right_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_7_Right_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_7_Right_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_7_Right_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_7_Right_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_7_Right_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_7_Right_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_7_Right_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_7_Right_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_7_Right_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_7_Right_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_7_Right_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_7_Right_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_7_Right_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_7_Right_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_7_Right_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_7_Right_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_7_Right_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_7_Right_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_7_Right_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_7_Right_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_7_Right_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_7_Right_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_7_Right_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_7_Right_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_7_Right_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_7_Right_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_7_Right_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_7_Right_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_7_Right_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_7_Right_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_7_Right_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_7_Right_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_7_Right_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_7_Right_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_8_Left_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_8_Left_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_8_Left_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_8_Left_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_8_Left_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_8_Left_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_8_Left_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_8_Left_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_8_Left_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_8_Left_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_8_Left_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_8_Left_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_8_Left_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_8_Left_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_8_Left_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_8_Left_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_8_Left_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_8_Left_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_8_Left_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_8_Left_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_8_Left_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_8_Left_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_8_Left_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_8_Left_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_8_Left_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_8_Left_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_8_Left_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_8_Left_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_8_Left_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_8_Left_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_8_Left_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_8_Left_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_8_Left_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_8_Left_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_8_Left_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_8_Left_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_8_Left_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_8_Left_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_8_Left_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_8_Left_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_8_Left_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_8_Left_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_8_Left_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_8_Left_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_8_Left_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_8_Left_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_8_Left_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_8_Left_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_8_Left_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_8_Left_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_8_Left_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_8_Left_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_8_Left_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_8_Left_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_8_Left_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_8_Left_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_8_Left_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_8_Left_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_8_Left_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_8_Left_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_8_Left_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_8_Left_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_8_Left_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_8_Left_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_8_Left_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_8_Left_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_8_Left_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_8_Left_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_8_Left_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_8_Left_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_8_Left_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_8_Left_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_8_Left_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_8_Left_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_8_Left_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_8_Left_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_8_Left_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_8_Left_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_8_Left_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_8_Left_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_8_Left_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_8_Left_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_8_Left_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_8_Left_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_8_Left_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_8_Left_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_8_Left_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_8_Left_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_8_Left_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_8_Left_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_8_Left_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_8_Left_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_8_Left_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_8_Left_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_8_Left_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_8_Left_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_8_Left_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_8_Left_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_8_Left_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_8_Left_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_8_Left_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_8_Left_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_8_Left_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_8_Left_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_8_Left_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_8_Left_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_8_Left_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_8_Left_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_8_Left_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_8_Left_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_8_Left_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_8_Left_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_8_Left_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_8_Left_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_8_Left_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_8_Left_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_8_Left_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_8_Left_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_8_Left_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_8_Left_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_8_Left_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_8_Left_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_8_Left_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_8_Left_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_8_Left_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_8_Left_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_8_Left_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_8_Left_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_8_Left_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_8_Left_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_8_Left_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_8_Left_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_8_Left_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_8_Left_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_8_Left_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_8_Left_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_8_Left_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_8_Left_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_8_Left_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_8_Left_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_8_Left_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_8_Left_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_8_Left_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_8_Left_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_8_Left_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_8_Left_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_8_Left_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_8_Left_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_8_Left_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_8_Left_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_8_Left_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_8_Left_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_8_Left_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_8_Left_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_8_Left_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_8_Left_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_8_Left_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_8_Left_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_8_Left_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_8_Left_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_8_Left_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_8_Left_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_8_Left_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_8_Left_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_8_Left_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_8_Left_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_8_Left_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_8_Left_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_8_Left_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_8_Left_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_8_Left_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_8_Left_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_8_Left_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_8_Left_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_8_Left_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_8_Left_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_8_Left_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_8_Left_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_8_Left_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_8_Left_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_8_Left_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_8_Left_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_8_Left_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_8_Left_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_8_Left_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_8_Left_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_8_Left_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_8_Left_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_8_Left_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_8_Left_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_8_Left_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_8_Left_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_8_Left_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_8_Left_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_8_Left_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_8_Left_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_8_Left_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_8_Left_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_8_Left_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_8_Left_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_8_Left_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_8_Left_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_8_Left_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_8_Left_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_8_Left_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_8_Left_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_8_Left_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_8_Left_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_8_Left_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_8_Left_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_8_Left_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_8_Left_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_8_Left_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_8_Left_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_8_Left_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_8_Left_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_8_Left_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_8_Left_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_8_Left_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_8_Left_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_8_Left_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_8_Left_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_8_Left_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_8_Left_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_8_Left_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_8_Left_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_8_Left_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_8_Left_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_8_Left_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_8_Left_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_8_Left_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_8_Left_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_8_Left_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_8_Left_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_8_Left_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_8_Left_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_8_Left_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_8_Left_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_8_Left_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_8_Left_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_8_Left_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_8_Left_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_8_Left_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_8_Left_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_8_Left_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_8_Left_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_8_Left_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_8_Left_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_8_Left_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_8_Left_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_8_Left_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_8_Left_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_8_Left_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_8_Left_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_8_Left_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_8_Left_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_8_Left_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_8_Left_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_8_Left_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_8_Left_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_8_Left_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_8_Left_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_8_Left_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_8_Left_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_8_Left_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_8_Left_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_8_Left_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_8_Left_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_8_Left_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_8_Left_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_8_Left_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_8_Left_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_8_Left_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_8_Left_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_8_Left_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_8_Left_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_8_Left_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_8_Left_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_8_Left_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_8_Left_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_8_Left_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_8_Left_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_8_Left_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_8_Left_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_8_Left_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_8_Left_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_8_Left_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_8_Left_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_8_Left_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_8_Left_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_8_Left_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_8_Left_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_8_Left_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_8_Left_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_8_Left_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_8_Left_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_8_Left_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_8_Left_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_8_Left_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_8_Left_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_8_Left_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_8_Left_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_8_Left_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_8_Left_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_8_Left_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_8_Left_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_8_Left_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_8_Left_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_8_Left_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_8_Left_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_8_Left_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_8_Left_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_8_Left_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_8_Left_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_8_Left_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_8_Left_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_8_Left_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_8_Left_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_8_Left_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_8_Left_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_8_Left_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_8_Left_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_8_Left_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_8_Left_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_8_Right_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_8_Right_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_8_Right_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_8_Right_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_8_Right_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_8_Right_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_8_Right_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_8_Right_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_8_Right_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_8_Right_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_8_Right_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_8_Right_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_8_Right_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_8_Right_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_8_Right_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_8_Right_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_8_Right_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_8_Right_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_8_Right_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_8_Right_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_8_Right_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_8_Right_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_8_Right_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_8_Right_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_8_Right_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_8_Right_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_8_Right_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_8_Right_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_8_Right_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_8_Right_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_8_Right_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_8_Right_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_8_Right_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_8_Right_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_8_Right_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_8_Right_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_8_Right_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_8_Right_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_8_Right_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_8_Right_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_8_Right_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_8_Right_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_8_Right_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_8_Right_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_8_Right_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_8_Right_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_8_Right_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_8_Right_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_8_Right_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_8_Right_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_8_Right_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_8_Right_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_8_Right_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_8_Right_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_8_Right_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_8_Right_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_8_Right_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_8_Right_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_8_Right_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_8_Right_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_8_Right_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_8_Right_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_8_Right_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_8_Right_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_8_Right_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_8_Right_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_8_Right_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_8_Right_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_8_Right_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_8_Right_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_8_Right_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_8_Right_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_8_Right_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_8_Right_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_8_Right_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_8_Right_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_8_Right_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_8_Right_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_8_Right_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_8_Right_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_8_Right_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_8_Right_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_8_Right_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_8_Right_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_8_Right_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_8_Right_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_8_Right_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_8_Right_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_8_Right_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_8_Right_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_8_Right_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_8_Right_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_8_Right_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_8_Right_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_8_Right_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_8_Right_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_8_Right_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_8_Right_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_8_Right_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_8_Right_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_8_Right_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_8_Right_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_8_Right_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_8_Right_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_8_Right_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_8_Right_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_8_Right_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_8_Right_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_8_Right_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_8_Right_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_8_Right_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_8_Right_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_8_Right_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_8_Right_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_8_Right_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_8_Right_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_8_Right_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_8_Right_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_8_Right_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_8_Right_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_8_Right_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_8_Right_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_8_Right_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_8_Right_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_8_Right_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_8_Right_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_8_Right_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_8_Right_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_8_Right_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_8_Right_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_8_Right_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_8_Right_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_8_Right_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_8_Right_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_8_Right_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_8_Right_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_8_Right_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_8_Right_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_8_Right_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_8_Right_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_8_Right_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_8_Right_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_8_Right_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_8_Right_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_8_Right_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_8_Right_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_8_Right_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_8_Right_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_8_Right_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_8_Right_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_8_Right_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_8_Right_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_8_Right_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_8_Right_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_8_Right_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_8_Right_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_8_Right_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_8_Right_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_8_Right_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_8_Right_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_8_Right_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_8_Right_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_8_Right_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_8_Right_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_8_Right_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_8_Right_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_8_Right_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_8_Right_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_8_Right_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_8_Right_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_8_Right_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_8_Right_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_8_Right_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_8_Right_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_8_Right_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_8_Right_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_8_Right_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_8_Right_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_8_Right_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_8_Right_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_8_Right_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_8_Right_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_8_Right_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_8_Right_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_8_Right_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_8_Right_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_8_Right_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_8_Right_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_8_Right_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_8_Right_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_8_Right_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_8_Right_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_8_Right_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_8_Right_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_8_Right_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_8_Right_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_8_Right_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_8_Right_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_8_Right_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_8_Right_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_8_Right_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_8_Right_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_8_Right_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_8_Right_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_8_Right_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_8_Right_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_8_Right_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_8_Right_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_8_Right_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_8_Right_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_8_Right_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_8_Right_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_8_Right_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_8_Right_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_8_Right_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_8_Right_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_8_Right_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_8_Right_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_8_Right_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_8_Right_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_8_Right_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_8_Right_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_8_Right_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_8_Right_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_8_Right_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_8_Right_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_8_Right_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_8_Right_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_8_Right_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_8_Right_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_8_Right_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_8_Right_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_8_Right_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_8_Right_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_8_Right_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_8_Right_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_8_Right_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_8_Right_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_8_Right_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_8_Right_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_8_Right_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_8_Right_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_8_Right_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_8_Right_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_8_Right_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_8_Right_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_8_Right_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_8_Right_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_8_Right_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_8_Right_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_8_Right_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_8_Right_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_8_Right_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_8_Right_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_8_Right_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_8_Right_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_8_Right_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_8_Right_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_8_Right_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_8_Right_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_8_Right_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_8_Right_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_8_Right_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_8_Right_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_8_Right_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_8_Right_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_8_Right_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_8_Right_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_8_Right_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_8_Right_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_8_Right_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_8_Right_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_8_Right_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_8_Right_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_8_Right_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_8_Right_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_8_Right_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_8_Right_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_8_Right_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_8_Right_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_8_Right_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_8_Right_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_8_Right_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_8_Right_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_8_Right_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_8_Right_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_8_Right_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_8_Right_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_8_Right_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_8_Right_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_8_Right_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_8_Right_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_8_Right_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_8_Right_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_8_Right_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_8_Right_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_8_Right_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_8_Right_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_8_Right_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_8_Right_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_8_Right_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_8_Right_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_8_Right_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_8_Right_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_8_Right_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_8_Right_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_8_Right_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_8_Right_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_8_Right_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_8_Right_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_8_Right_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_8_Right_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_8_Right_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_8_Right_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_8_Right_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_8_Right_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_8_Right_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_8_Right_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_8_Right_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_8_Right_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_8_Right_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_8_Right_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_8_Right_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_8_Right_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_9_Left_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_9_Left_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_9_Left_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_9_Left_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_9_Left_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_9_Left_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_9_Left_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_9_Left_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_9_Left_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_9_Left_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_9_Left_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_9_Left_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_9_Left_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_9_Left_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_9_Left_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_9_Left_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_9_Left_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_9_Left_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_9_Left_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_9_Left_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_9_Left_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_9_Left_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_9_Left_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_9_Left_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_9_Left_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_9_Left_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_9_Left_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_9_Left_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_9_Left_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_9_Left_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_9_Left_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_9_Left_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_9_Left_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_9_Left_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_9_Left_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_9_Left_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_9_Left_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_9_Left_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_9_Left_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_9_Left_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_9_Left_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_9_Left_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_9_Left_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_9_Left_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_9_Left_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_9_Left_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_9_Left_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_9_Left_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_9_Left_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_9_Left_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_9_Left_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_9_Left_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_9_Left_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_9_Left_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_9_Left_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_9_Left_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_9_Left_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_9_Left_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_9_Left_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_9_Left_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_9_Left_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_9_Left_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_9_Left_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_9_Left_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_9_Left_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_9_Left_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_9_Left_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_9_Left_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_9_Left_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_9_Left_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_9_Left_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_9_Left_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_9_Left_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_9_Left_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_9_Left_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_9_Left_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_9_Left_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_9_Left_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_9_Left_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_9_Left_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_9_Left_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_9_Left_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_9_Left_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_9_Left_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_9_Left_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_9_Left_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_9_Left_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_9_Left_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_9_Left_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_9_Left_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_9_Left_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_9_Left_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_9_Left_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_9_Left_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_9_Left_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_9_Left_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_9_Left_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_9_Left_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_9_Left_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_9_Left_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_9_Left_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_9_Left_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_9_Left_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_9_Left_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_9_Left_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_9_Left_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_9_Left_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_9_Left_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_9_Left_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_9_Left_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_9_Left_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_9_Left_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_9_Left_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_9_Left_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_9_Left_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_9_Left_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_9_Left_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_9_Left_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_9_Left_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_9_Left_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_9_Left_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_9_Left_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_9_Left_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_9_Left_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_9_Left_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_9_Left_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_9_Left_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_9_Left_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_9_Left_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_9_Left_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_9_Left_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_9_Left_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_9_Left_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_9_Left_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_9_Left_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_9_Left_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_9_Left_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_9_Left_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_9_Left_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_9_Left_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_9_Left_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_9_Left_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_9_Left_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_9_Left_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_9_Left_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_9_Left_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_9_Left_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_9_Left_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_9_Left_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_9_Left_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_9_Left_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_9_Left_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_9_Left_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_9_Left_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_9_Left_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_9_Left_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_9_Left_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_9_Left_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_9_Left_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_9_Left_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_9_Left_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_9_Left_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_9_Left_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_9_Left_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_9_Left_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_9_Left_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_9_Left_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_9_Left_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_9_Left_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_9_Left_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_9_Left_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_9_Left_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_9_Left_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_9_Left_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_9_Left_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_9_Left_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_9_Left_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_9_Left_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_9_Left_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_9_Left_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_9_Left_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_9_Left_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_9_Left_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_9_Left_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_9_Left_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_9_Left_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_9_Left_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_9_Left_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_9_Left_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_9_Left_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_9_Left_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_9_Left_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_9_Left_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_9_Left_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_9_Left_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_9_Left_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_9_Left_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_9_Left_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_9_Left_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_9_Left_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_9_Left_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_9_Left_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_9_Left_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_9_Left_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_9_Left_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_9_Left_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_9_Left_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_9_Left_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_9_Left_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_9_Left_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_9_Left_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_9_Left_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_9_Left_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_9_Left_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_9_Left_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_9_Left_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_9_Left_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_9_Left_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_9_Left_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_9_Left_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_9_Left_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_9_Left_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_9_Left_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_9_Left_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_9_Left_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_9_Left_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_9_Left_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_9_Left_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_9_Left_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_9_Left_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_9_Left_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_9_Left_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_9_Left_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_9_Left_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_9_Left_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_9_Left_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_9_Left_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_9_Left_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_9_Left_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_9_Left_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_9_Left_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_9_Left_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_9_Left_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_9_Left_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_9_Left_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_9_Left_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_9_Left_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_9_Left_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_9_Left_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_9_Left_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_9_Left_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_9_Left_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_9_Left_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_9_Left_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_9_Left_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_9_Left_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_9_Left_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_9_Left_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_9_Left_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_9_Left_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_9_Left_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_9_Left_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_9_Left_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_9_Left_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_9_Left_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_9_Left_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_9_Left_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_9_Left_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_9_Left_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_9_Left_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_9_Left_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_9_Left_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_9_Left_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_9_Left_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_9_Left_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_9_Left_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_9_Left_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_9_Left_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_9_Left_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_9_Left_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_9_Left_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_9_Left_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_9_Left_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_9_Left_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_9_Left_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_9_Left_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_9_Left_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_9_Left_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_9_Left_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_9_Left_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_9_Left_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_9_Left_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_9_Left_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_9_Left_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_9_Left_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_9_Left_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_9_Left_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_9_Left_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_9_Left_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_9_Left_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_9_Left_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_9_Left_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_9_Left_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_9_Left_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_9_Left_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_9_Left_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_9_Left_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_9_Left_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_9_Left_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_9_Left_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_9_Left_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_9_Left_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_9_Left_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_9_Left_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_9_Left_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_9_Left_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_9_Left_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_9_Left_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_9_Left_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_9_Left_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_9_Left_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_9_Left_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_9_Left_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_9_Left_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_9_Right_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_9_Right_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_9_Right_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_9_Right_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_9_Right_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_9_Right_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_9_Right_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_9_Right_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_9_Right_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_9_Right_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_9_Right_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_9_Right_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_9_Right_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_9_Right_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_9_Right_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_9_Right_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_9_Right_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_9_Right_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_9_Right_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_9_Right_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_9_Right_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_9_Right_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_9_Right_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_9_Right_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_9_Right_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_9_Right_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_9_Right_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_9_Right_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_9_Right_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_9_Right_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_9_Right_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_9_Right_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_9_Right_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_9_Right_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_9_Right_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_9_Right_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_9_Right_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_9_Right_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_9_Right_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_9_Right_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_9_Right_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_9_Right_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_9_Right_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_9_Right_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_9_Right_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_9_Right_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_9_Right_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_9_Right_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_9_Right_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_9_Right_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_9_Right_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_9_Right_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_9_Right_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_9_Right_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_9_Right_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_9_Right_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_9_Right_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_9_Right_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_9_Right_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_9_Right_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_9_Right_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_9_Right_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_9_Right_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_9_Right_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_9_Right_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_9_Right_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_9_Right_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_9_Right_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_9_Right_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_9_Right_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_9_Right_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_9_Right_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_9_Right_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_9_Right_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_9_Right_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_9_Right_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_9_Right_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_9_Right_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_9_Right_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_9_Right_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_9_Right_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_9_Right_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_9_Right_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_9_Right_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_9_Right_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_9_Right_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_9_Right_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_9_Right_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_9_Right_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_9_Right_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_9_Right_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_9_Right_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_9_Right_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_9_Right_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_9_Right_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_9_Right_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_9_Right_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_9_Right_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_9_Right_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_9_Right_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_9_Right_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_9_Right_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_9_Right_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_9_Right_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_9_Right_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_9_Right_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_9_Right_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_9_Right_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_9_Right_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_9_Right_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_9_Right_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_9_Right_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_9_Right_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_9_Right_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_9_Right_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_9_Right_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_9_Right_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_9_Right_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_9_Right_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_9_Right_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_9_Right_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_9_Right_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_9_Right_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_9_Right_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_9_Right_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_9_Right_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_9_Right_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_9_Right_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_9_Right_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_9_Right_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_9_Right_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_9_Right_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_9_Right_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_9_Right_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_9_Right_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_9_Right_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_9_Right_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_9_Right_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_9_Right_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_9_Right_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_9_Right_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_9_Right_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_9_Right_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_9_Right_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_9_Right_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_9_Right_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_9_Right_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_9_Right_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_9_Right_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_9_Right_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_9_Right_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_9_Right_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_9_Right_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_9_Right_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_9_Right_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_9_Right_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_9_Right_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_9_Right_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_9_Right_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_9_Right_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_9_Right_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_9_Right_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_9_Right_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_9_Right_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_9_Right_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_9_Right_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_9_Right_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_9_Right_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_9_Right_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_9_Right_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_9_Right_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_9_Right_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_9_Right_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_9_Right_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_9_Right_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_9_Right_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_9_Right_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_9_Right_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_9_Right_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_9_Right_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_9_Right_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_9_Right_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_9_Right_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_9_Right_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_9_Right_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_9_Right_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_9_Right_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_9_Right_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_9_Right_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_9_Right_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_9_Right_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_9_Right_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_9_Right_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_9_Right_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_9_Right_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_9_Right_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_9_Right_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_9_Right_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_9_Right_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_9_Right_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_9_Right_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_9_Right_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_9_Right_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_9_Right_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_9_Right_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_9_Right_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_9_Right_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_9_Right_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_9_Right_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_9_Right_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_9_Right_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_9_Right_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_9_Right_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_9_Right_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_9_Right_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_9_Right_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_9_Right_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_9_Right_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_9_Right_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_9_Right_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_9_Right_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_9_Right_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_9_Right_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_9_Right_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_9_Right_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_9_Right_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_9_Right_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_9_Right_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_9_Right_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_9_Right_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_9_Right_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_9_Right_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_9_Right_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_9_Right_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_9_Right_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_9_Right_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_9_Right_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_9_Right_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_9_Right_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_9_Right_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_9_Right_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_9_Right_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_9_Right_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_9_Right_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_9_Right_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_9_Right_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_9_Right_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_9_Right_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_9_Right_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_9_Right_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_9_Right_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_9_Right_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_9_Right_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_9_Right_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_9_Right_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_9_Right_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_9_Right_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_9_Right_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_9_Right_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_9_Right_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_9_Right_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_9_Right_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_9_Right_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_9_Right_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_9_Right_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_9_Right_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_9_Right_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_9_Right_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_9_Right_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_9_Right_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_9_Right_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_9_Right_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_9_Right_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_9_Right_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_9_Right_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_9_Right_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_9_Right_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_9_Right_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_9_Right_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_9_Right_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_9_Right_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_9_Right_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_9_Right_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_9_Right_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_9_Right_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_9_Right_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_9_Right_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_9_Right_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_9_Right_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_9_Right_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_9_Right_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_9_Right_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_9_Right_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_9_Right_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_9_Right_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_9_Right_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_9_Right_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_9_Right_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_9_Right_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_9_Right_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_9_Right_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_9_Right_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_9_Right_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_9_Right_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_9_Right_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_9_Right_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_9_Right_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_9_Right_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_9_Right_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_9_Right_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_9_Right_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_9_Right_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_9_Right_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_9_Right_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_9_Right_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_9_Right_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_9_Right_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_9_Right_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_9_Right_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_9_Right_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_9_Right_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_9_Right_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_9_Right_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_9_Right_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_10_Left_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_10_Left_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_10_Left_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_10_Left_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_10_Left_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_10_Left_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_10_Left_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_10_Left_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_10_Left_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_10_Left_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_10_Left_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_10_Left_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_10_Left_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_10_Left_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_10_Left_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_10_Left_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_10_Left_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_10_Left_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_10_Left_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_10_Left_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_10_Left_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_10_Left_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_10_Left_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_10_Left_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_10_Left_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_10_Left_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_10_Left_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_10_Left_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_10_Left_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_10_Left_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_10_Left_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_10_Left_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_10_Left_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_10_Left_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_10_Left_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_10_Left_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_10_Left_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_10_Left_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_10_Left_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_10_Left_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_10_Left_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_10_Left_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_10_Left_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_10_Left_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_10_Left_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_10_Left_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_10_Left_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_10_Left_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_10_Left_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_10_Left_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_10_Left_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_10_Left_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_10_Left_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_10_Left_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_10_Left_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_10_Left_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_10_Left_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_10_Left_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_10_Left_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_10_Left_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_10_Left_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_10_Left_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_10_Left_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_10_Left_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_10_Left_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_10_Left_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_10_Left_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_10_Left_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_10_Left_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_10_Left_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_10_Left_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_10_Left_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_10_Left_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_10_Left_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_10_Left_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_10_Left_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_10_Left_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_10_Left_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_10_Left_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_10_Left_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_10_Left_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_10_Left_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_10_Left_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_10_Left_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_10_Left_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_10_Left_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_10_Left_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_10_Left_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_10_Left_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_10_Left_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_10_Left_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_10_Left_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_10_Left_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_10_Left_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_10_Left_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_10_Left_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_10_Left_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_10_Left_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_10_Left_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_10_Left_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_10_Left_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_10_Left_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_10_Left_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_10_Left_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_10_Left_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_10_Left_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_10_Left_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_10_Left_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_10_Left_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_10_Left_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_10_Left_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_10_Left_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_10_Left_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_10_Left_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_10_Left_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_10_Left_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_10_Left_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_10_Left_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_10_Left_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_10_Left_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_10_Left_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_10_Left_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_10_Left_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_10_Left_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_10_Left_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_10_Left_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_10_Left_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_10_Left_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_10_Left_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_10_Left_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_10_Left_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_10_Left_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_10_Left_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_10_Left_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_10_Left_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_10_Left_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_10_Left_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_10_Left_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_10_Left_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_10_Left_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_10_Left_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_10_Left_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_10_Left_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_10_Left_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_10_Left_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_10_Left_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_10_Left_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_10_Left_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_10_Left_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_10_Left_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_10_Left_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_10_Left_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_10_Left_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_10_Left_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_10_Left_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_10_Left_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_10_Left_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_10_Left_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_10_Left_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_10_Left_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_10_Left_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_10_Left_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_10_Left_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_10_Left_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_10_Left_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_10_Left_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_10_Left_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_10_Left_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_10_Left_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_10_Left_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_10_Left_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_10_Left_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_10_Left_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_10_Left_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_10_Left_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_10_Left_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_10_Left_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_10_Left_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_10_Left_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_10_Left_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_10_Left_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_10_Left_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_10_Left_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_10_Left_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_10_Left_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_10_Left_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_10_Left_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_10_Left_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_10_Left_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_10_Left_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_10_Left_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_10_Left_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_10_Left_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_10_Left_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_10_Left_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_10_Left_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_10_Left_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_10_Left_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_10_Left_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_10_Left_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_10_Left_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_10_Left_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_10_Left_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_10_Left_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_10_Left_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_10_Left_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_10_Left_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_10_Left_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_10_Left_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_10_Left_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_10_Left_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_10_Left_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_10_Left_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_10_Left_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_10_Left_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_10_Left_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_10_Left_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_10_Left_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_10_Left_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_10_Left_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_10_Left_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_10_Left_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_10_Left_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_10_Left_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_10_Left_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_10_Left_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_10_Left_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_10_Left_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_10_Left_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_10_Left_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_10_Left_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_10_Left_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_10_Left_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_10_Left_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_10_Left_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_10_Left_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_10_Left_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_10_Left_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_10_Left_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_10_Left_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_10_Left_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_10_Left_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_10_Left_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_10_Left_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_10_Left_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_10_Left_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_10_Left_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_10_Left_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_10_Left_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_10_Left_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_10_Left_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_10_Left_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_10_Left_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_10_Left_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_10_Left_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_10_Left_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_10_Left_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_10_Left_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_10_Left_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_10_Left_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_10_Left_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_10_Left_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_10_Left_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_10_Left_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_10_Left_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_10_Left_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_10_Left_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_10_Left_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_10_Left_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_10_Left_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_10_Left_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_10_Left_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_10_Left_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_10_Left_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_10_Left_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_10_Left_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_10_Left_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_10_Left_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_10_Left_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_10_Left_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_10_Left_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_10_Left_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_10_Left_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_10_Left_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_10_Left_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_10_Left_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_10_Left_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_10_Left_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_10_Left_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_10_Left_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_10_Left_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_10_Left_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_10_Left_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_10_Left_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_10_Left_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_10_Left_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_10_Left_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_10_Left_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_10_Left_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_10_Left_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_10_Left_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_10_Left_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_10_Left_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_10_Left_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_10_Left_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_10_Left_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_10_Left_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_10_Left_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_10_Left_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_10_Left_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_10_Left_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_10_Left_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_10_Left_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_10_Left_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_10_Left_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_10_Left_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_10_Left_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_10_Left_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_10_Left_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_10_Left_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_10_Left_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_10_Left_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_10_Left_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_10_Left_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_10_Right_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_10_Right_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_10_Right_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_10_Right_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_10_Right_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_10_Right_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_10_Right_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_10_Right_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_10_Right_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_10_Right_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_10_Right_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_10_Right_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_10_Right_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_10_Right_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_10_Right_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_10_Right_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_10_Right_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_10_Right_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_10_Right_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_10_Right_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_10_Right_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_10_Right_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_10_Right_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_10_Right_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_10_Right_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_10_Right_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_10_Right_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_10_Right_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_10_Right_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_10_Right_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_10_Right_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_10_Right_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_10_Right_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_10_Right_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_10_Right_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_10_Right_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_10_Right_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_10_Right_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_10_Right_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_10_Right_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_10_Right_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_10_Right_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_10_Right_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_10_Right_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_10_Right_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_10_Right_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_10_Right_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_10_Right_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_10_Right_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_10_Right_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_10_Right_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_10_Right_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_10_Right_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_10_Right_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_10_Right_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_10_Right_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_10_Right_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_10_Right_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_10_Right_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_10_Right_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_10_Right_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_10_Right_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_10_Right_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_10_Right_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_10_Right_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_10_Right_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_10_Right_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_10_Right_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_10_Right_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_10_Right_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_10_Right_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_10_Right_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_10_Right_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_10_Right_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_10_Right_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_10_Right_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_10_Right_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_10_Right_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_10_Right_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_10_Right_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_10_Right_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_10_Right_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_10_Right_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_10_Right_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_10_Right_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_10_Right_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_10_Right_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_10_Right_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_10_Right_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_10_Right_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_10_Right_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_10_Right_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_10_Right_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_10_Right_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_10_Right_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_10_Right_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_10_Right_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_10_Right_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_10_Right_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_10_Right_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_10_Right_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_10_Right_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_10_Right_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_10_Right_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_10_Right_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_10_Right_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_10_Right_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_10_Right_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_10_Right_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_10_Right_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_10_Right_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_10_Right_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_10_Right_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_10_Right_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_10_Right_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_10_Right_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_10_Right_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_10_Right_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_10_Right_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_10_Right_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_10_Right_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_10_Right_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_10_Right_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_10_Right_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_10_Right_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_10_Right_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_10_Right_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_10_Right_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_10_Right_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_10_Right_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_10_Right_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_10_Right_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_10_Right_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_10_Right_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_10_Right_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_10_Right_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_10_Right_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_10_Right_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_10_Right_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_10_Right_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_10_Right_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_10_Right_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_10_Right_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_10_Right_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_10_Right_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_10_Right_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_10_Right_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_10_Right_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_10_Right_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_10_Right_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_10_Right_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_10_Right_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_10_Right_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_10_Right_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_10_Right_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_10_Right_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_10_Right_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_10_Right_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_10_Right_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_10_Right_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_10_Right_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_10_Right_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_10_Right_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_10_Right_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_10_Right_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_10_Right_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_10_Right_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_10_Right_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_10_Right_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_10_Right_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_10_Right_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_10_Right_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_10_Right_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_10_Right_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_10_Right_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_10_Right_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_10_Right_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_10_Right_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_10_Right_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_10_Right_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_10_Right_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_10_Right_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_10_Right_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_10_Right_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_10_Right_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_10_Right_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_10_Right_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_10_Right_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_10_Right_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_10_Right_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_10_Right_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_10_Right_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_10_Right_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_10_Right_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_10_Right_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_10_Right_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_10_Right_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_10_Right_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_10_Right_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_10_Right_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_10_Right_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_10_Right_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_10_Right_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_10_Right_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_10_Right_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_10_Right_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_10_Right_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_10_Right_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_10_Right_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_10_Right_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_10_Right_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_10_Right_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_10_Right_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_10_Right_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_10_Right_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_10_Right_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_10_Right_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_10_Right_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_10_Right_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_10_Right_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_10_Right_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_10_Right_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_10_Right_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_10_Right_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_10_Right_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_10_Right_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_10_Right_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_10_Right_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_10_Right_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_10_Right_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_10_Right_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_10_Right_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_10_Right_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_10_Right_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_10_Right_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_10_Right_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_10_Right_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_10_Right_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_10_Right_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_10_Right_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_10_Right_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_10_Right_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_10_Right_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_10_Right_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_10_Right_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_10_Right_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_10_Right_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_10_Right_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_10_Right_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_10_Right_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_10_Right_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_10_Right_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_10_Right_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_10_Right_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_10_Right_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_10_Right_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_10_Right_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_10_Right_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_10_Right_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_10_Right_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_10_Right_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_10_Right_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_10_Right_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_10_Right_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_10_Right_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_10_Right_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_10_Right_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_10_Right_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_10_Right_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_10_Right_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_10_Right_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_10_Right_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_10_Right_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_10_Right_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_10_Right_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_10_Right_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_10_Right_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_10_Right_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_10_Right_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_10_Right_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_10_Right_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_10_Right_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_10_Right_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_10_Right_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_10_Right_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_10_Right_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_10_Right_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_10_Right_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_10_Right_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_10_Right_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_10_Right_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_10_Right_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_10_Right_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_10_Right_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_10_Right_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_10_Right_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_10_Right_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_10_Right_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_10_Right_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_10_Right_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_10_Right_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_10_Right_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_10_Right_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_10_Right_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_10_Right_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_10_Right_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_10_Right_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_10_Right_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_10_Right_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_10_Right_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_10_Right_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_10_Right_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_10_Right_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_10_Right_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_10_Right_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_10_Right_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_10_Right_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_10_Right_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_10_Right_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_10_Right_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_10_Right_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_10_Right_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_10_Right_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_10_Right_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_11_Left_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_11_Left_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_11_Left_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_11_Left_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_11_Left_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_11_Left_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_11_Left_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_11_Left_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_11_Left_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_11_Left_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_11_Left_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_11_Left_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_11_Left_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_11_Left_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_11_Left_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_11_Left_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_11_Left_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_11_Left_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_11_Left_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_11_Left_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_11_Left_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_11_Left_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_11_Left_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_11_Left_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_11_Left_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_11_Left_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_11_Left_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_11_Left_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_11_Left_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_11_Left_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_11_Left_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_11_Left_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_11_Left_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_11_Left_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_11_Left_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_11_Left_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_11_Left_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_11_Left_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_11_Left_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_11_Left_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_11_Left_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_11_Left_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_11_Left_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_11_Left_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_11_Left_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_11_Left_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_11_Left_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_11_Left_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_11_Left_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_11_Left_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_11_Left_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_11_Left_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_11_Left_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_11_Left_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_11_Left_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_11_Left_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_11_Left_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_11_Left_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_11_Left_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_11_Left_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_11_Left_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_11_Left_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_11_Left_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_11_Left_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_11_Left_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_11_Left_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_11_Left_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_11_Left_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_11_Left_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_11_Left_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_11_Left_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_11_Left_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_11_Left_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_11_Left_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_11_Left_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_11_Left_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_11_Left_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_11_Left_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_11_Left_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_11_Left_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_11_Left_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_11_Left_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_11_Left_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_11_Left_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_11_Left_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_11_Left_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_11_Left_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_11_Left_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_11_Left_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_11_Left_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_11_Left_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_11_Left_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_11_Left_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_11_Left_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_11_Left_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_11_Left_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_11_Left_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_11_Left_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_11_Left_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_11_Left_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_11_Left_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_11_Left_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_11_Left_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_11_Left_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_11_Left_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_11_Left_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_11_Left_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_11_Left_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_11_Left_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_11_Left_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_11_Left_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_11_Left_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_11_Left_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_11_Left_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_11_Left_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_11_Left_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_11_Left_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_11_Left_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_11_Left_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_11_Left_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_11_Left_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_11_Left_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_11_Left_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_11_Left_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_11_Left_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_11_Left_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_11_Left_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_11_Left_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_11_Left_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_11_Left_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_11_Left_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_11_Left_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_11_Left_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_11_Left_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_11_Left_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_11_Left_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_11_Left_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_11_Left_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_11_Left_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_11_Left_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_11_Left_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_11_Left_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_11_Left_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_11_Left_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_11_Left_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_11_Left_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_11_Left_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_11_Left_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_11_Left_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_11_Left_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_11_Left_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_11_Left_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_11_Left_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_11_Left_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_11_Left_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_11_Left_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_11_Left_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_11_Left_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_11_Left_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_11_Left_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_11_Left_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_11_Left_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_11_Left_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_11_Left_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_11_Left_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_11_Left_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_11_Left_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_11_Left_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_11_Left_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_11_Left_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_11_Left_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_11_Left_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_11_Left_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_11_Left_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_11_Left_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_11_Left_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_11_Left_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_11_Left_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_11_Left_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_11_Left_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_11_Left_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_11_Left_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_11_Left_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_11_Left_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_11_Left_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_11_Left_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_11_Left_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_11_Left_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_11_Left_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_11_Left_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_11_Left_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_11_Left_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_11_Left_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_11_Left_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_11_Left_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_11_Left_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_11_Left_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_11_Left_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_11_Left_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_11_Left_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_11_Left_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_11_Left_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_11_Left_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_11_Left_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_11_Left_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_11_Left_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_11_Left_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_11_Left_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_11_Left_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_11_Left_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_11_Left_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_11_Left_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_11_Left_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_11_Left_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_11_Left_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_11_Left_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_11_Left_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_11_Left_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_11_Left_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_11_Left_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_11_Left_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_11_Left_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_11_Left_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_11_Left_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_11_Left_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_11_Left_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_11_Left_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_11_Left_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_11_Left_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_11_Left_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_11_Left_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_11_Left_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_11_Left_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_11_Left_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_11_Left_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_11_Left_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_11_Left_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_11_Left_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_11_Left_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_11_Left_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_11_Left_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_11_Left_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_11_Left_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_11_Left_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_11_Left_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_11_Left_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_11_Left_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_11_Left_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_11_Left_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_11_Left_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_11_Left_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_11_Left_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_11_Left_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_11_Left_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_11_Left_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_11_Left_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_11_Left_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_11_Left_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_11_Left_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_11_Left_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_11_Left_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_11_Left_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_11_Left_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_11_Left_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_11_Left_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_11_Left_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_11_Left_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_11_Left_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_11_Left_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_11_Left_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_11_Left_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_11_Left_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_11_Left_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_11_Left_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_11_Left_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_11_Left_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_11_Left_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_11_Left_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_11_Left_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_11_Left_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_11_Left_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_11_Left_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_11_Left_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_11_Left_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_11_Left_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_11_Left_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_11_Left_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_11_Left_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_11_Left_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_11_Left_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_11_Left_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_11_Left_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_11_Left_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_11_Left_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_11_Left_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_11_Left_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_11_Left_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_11_Left_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_11_Left_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_11_Left_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_11_Left_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_11_Left_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_11_Left_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_11_Left_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_11_Left_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_11_Left_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_11_Left_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_11_Left_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_11_Left_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_11_Left_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_11_Left_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_11_Left_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_11_Left_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_11_Left_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_11_Left_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_11_Left_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_11_Left_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_11_Left_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_11_Left_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_11_Left_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_11_Left_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_11_Left_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_11_Left_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_11_Left_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_11_Right_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_11_Right_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_11_Right_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_11_Right_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_11_Right_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_11_Right_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_11_Right_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_11_Right_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_11_Right_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_11_Right_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_11_Right_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_11_Right_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_11_Right_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_11_Right_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_11_Right_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_11_Right_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_11_Right_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_11_Right_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_11_Right_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_11_Right_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_11_Right_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_11_Right_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_11_Right_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_11_Right_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_11_Right_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_11_Right_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_11_Right_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_11_Right_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_11_Right_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_11_Right_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_11_Right_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_11_Right_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_11_Right_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_11_Right_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_11_Right_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_11_Right_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_11_Right_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_11_Right_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_11_Right_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_11_Right_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_11_Right_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_11_Right_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_11_Right_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_11_Right_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_11_Right_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_11_Right_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_11_Right_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_11_Right_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_11_Right_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_11_Right_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_11_Right_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_11_Right_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_11_Right_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_11_Right_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_11_Right_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_11_Right_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_11_Right_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_11_Right_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_11_Right_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_11_Right_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_11_Right_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_11_Right_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_11_Right_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_11_Right_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_11_Right_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_11_Right_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_11_Right_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_11_Right_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_11_Right_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_11_Right_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_11_Right_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_11_Right_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_11_Right_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_11_Right_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_11_Right_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_11_Right_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_11_Right_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_11_Right_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_11_Right_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_11_Right_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_11_Right_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_11_Right_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_11_Right_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_11_Right_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_11_Right_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_11_Right_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_11_Right_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_11_Right_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_11_Right_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_11_Right_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_11_Right_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_11_Right_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_11_Right_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_11_Right_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_11_Right_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_11_Right_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_11_Right_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_11_Right_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_11_Right_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_11_Right_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_11_Right_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_11_Right_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_11_Right_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_11_Right_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_11_Right_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_11_Right_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_11_Right_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_11_Right_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_11_Right_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_11_Right_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_11_Right_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_11_Right_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_11_Right_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_11_Right_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_11_Right_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_11_Right_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_11_Right_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_11_Right_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_11_Right_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_11_Right_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_11_Right_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_11_Right_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_11_Right_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_11_Right_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_11_Right_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_11_Right_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_11_Right_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_11_Right_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_11_Right_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_11_Right_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_11_Right_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_11_Right_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_11_Right_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_11_Right_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_11_Right_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_11_Right_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_11_Right_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_11_Right_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_11_Right_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_11_Right_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_11_Right_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_11_Right_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_11_Right_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_11_Right_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_11_Right_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_11_Right_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_11_Right_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_11_Right_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_11_Right_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_11_Right_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_11_Right_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_11_Right_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_11_Right_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_11_Right_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_11_Right_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_11_Right_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_11_Right_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_11_Right_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_11_Right_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_11_Right_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_11_Right_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_11_Right_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_11_Right_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_11_Right_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_11_Right_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_11_Right_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_11_Right_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_11_Right_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_11_Right_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_11_Right_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_11_Right_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_11_Right_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_11_Right_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_11_Right_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_11_Right_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_11_Right_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_11_Right_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_11_Right_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_11_Right_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_11_Right_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_11_Right_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_11_Right_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_11_Right_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_11_Right_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_11_Right_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_11_Right_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_11_Right_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_11_Right_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_11_Right_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_11_Right_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_11_Right_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_11_Right_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_11_Right_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_11_Right_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_11_Right_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_11_Right_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_11_Right_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_11_Right_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_11_Right_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_11_Right_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_11_Right_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_11_Right_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_11_Right_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_11_Right_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_11_Right_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_11_Right_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_11_Right_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_11_Right_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_11_Right_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_11_Right_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_11_Right_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_11_Right_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_11_Right_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_11_Right_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_11_Right_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_11_Right_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_11_Right_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_11_Right_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_11_Right_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_11_Right_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_11_Right_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_11_Right_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_11_Right_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_11_Right_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_11_Right_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_11_Right_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_11_Right_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_11_Right_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_11_Right_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_11_Right_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_11_Right_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_11_Right_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_11_Right_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_11_Right_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_11_Right_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_11_Right_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_11_Right_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_11_Right_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_11_Right_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_11_Right_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_11_Right_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_11_Right_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_11_Right_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_11_Right_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_11_Right_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_11_Right_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_11_Right_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_11_Right_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_11_Right_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_11_Right_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_11_Right_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_11_Right_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_11_Right_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_11_Right_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_11_Right_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_11_Right_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_11_Right_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_11_Right_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_11_Right_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_11_Right_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_11_Right_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_11_Right_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_11_Right_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_11_Right_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_11_Right_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_11_Right_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_11_Right_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_11_Right_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_11_Right_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_11_Right_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_11_Right_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_11_Right_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_11_Right_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_11_Right_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_11_Right_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_11_Right_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_11_Right_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_11_Right_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_11_Right_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_11_Right_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_11_Right_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_11_Right_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_11_Right_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_11_Right_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_11_Right_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_11_Right_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_11_Right_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_11_Right_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_11_Right_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_11_Right_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_11_Right_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_11_Right_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_11_Right_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_11_Right_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_11_Right_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_11_Right_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_11_Right_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_11_Right_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_11_Right_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_11_Right_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_11_Right_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_11_Right_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_11_Right_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_11_Right_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_11_Right_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_11_Right_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_11_Right_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_11_Right_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_11_Right_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_11_Right_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_11_Right_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_11_Right_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_11_Right_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_11_Right_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_11_Right_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_11_Right_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_11_Right_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_11_Right_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_11_Right_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_11_Right_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_11_Right_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_11_Right_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_11_Right_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_11_Right_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_12_Left_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_12_Left_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_12_Left_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_12_Left_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_12_Left_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_12_Left_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_12_Left_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_12_Left_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_12_Left_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_12_Left_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_12_Left_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_12_Left_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_12_Left_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_12_Left_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_12_Left_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_12_Left_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_12_Left_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_12_Left_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_12_Left_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_12_Left_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_12_Left_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_12_Left_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_12_Left_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_12_Left_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_12_Left_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_12_Left_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_12_Left_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_12_Left_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_12_Left_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_12_Left_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_12_Left_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_12_Left_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_12_Left_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_12_Left_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_12_Left_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_12_Left_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_12_Left_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_12_Left_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_12_Left_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_12_Left_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_12_Left_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_12_Left_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_12_Left_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_12_Left_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_12_Left_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_12_Left_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_12_Left_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_12_Left_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_12_Left_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_12_Left_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_12_Left_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_12_Left_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_12_Left_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_12_Left_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_12_Left_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_12_Left_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_12_Left_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_12_Left_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_12_Left_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_12_Left_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_12_Left_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_12_Left_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_12_Left_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_12_Left_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_12_Left_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_12_Left_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_12_Left_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_12_Left_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_12_Left_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_12_Left_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_12_Left_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_12_Left_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_12_Left_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_12_Left_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_12_Left_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_12_Left_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_12_Left_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_12_Left_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_12_Left_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_12_Left_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_12_Left_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_12_Left_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_12_Left_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_12_Left_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_12_Left_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_12_Left_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_12_Left_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_12_Left_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_12_Left_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_12_Left_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_12_Left_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_12_Left_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_12_Left_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_12_Left_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_12_Left_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_12_Left_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_12_Left_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_12_Left_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_12_Left_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_12_Left_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_12_Left_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_12_Left_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_12_Left_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_12_Left_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_12_Left_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_12_Left_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_12_Left_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_12_Left_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_12_Left_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_12_Left_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_12_Left_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_12_Left_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_12_Left_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_12_Left_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_12_Left_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_12_Left_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_12_Left_6596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_12_Left_6597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_12_Left_6598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_12_Left_6599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_12_Left_6600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_12_Left_6601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_12_Left_6602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_12_Left_6603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_12_Left_6604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_12_Left_6605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_12_Left_6606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_12_Left_6607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_12_Left_6608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_12_Left_6609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_12_Left_6610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_12_Left_6611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_12_Left_6612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_12_Left_6613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_12_Left_6614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_12_Left_6615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_12_Left_6616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_12_Left_6617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_12_Left_6618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_12_Left_6619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_12_Left_6620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_12_Left_6621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_12_Left_6622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_12_Left_6623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_12_Left_6624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_12_Left_6625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_12_Left_6626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_12_Left_6627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_12_Left_6628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_12_Left_6629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_12_Left_6630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_12_Left_6631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_12_Left_6632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_12_Left_6633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_12_Left_6634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_12_Left_6635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_12_Left_6636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_12_Left_6637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_12_Left_6638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_12_Left_6639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_12_Left_6640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_12_Left_6641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_12_Left_6642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_12_Left_6643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_12_Left_6644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_12_Left_6645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_12_Left_6646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_12_Left_6647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_12_Left_6648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_12_Left_6649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_12_Left_6650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_12_Left_6651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_12_Left_6652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_12_Left_6653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_12_Left_6654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_12_Left_6655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_12_Left_6656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_12_Left_6657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_12_Left_6658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_12_Left_6659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_12_Left_6660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_12_Left_6661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_12_Left_6662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_12_Left_6663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_12_Left_6664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_12_Left_6665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_12_Left_6666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_12_Left_6667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_12_Left_6668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_12_Left_6669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_12_Left_6670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_12_Left_6671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_12_Left_6672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_12_Left_6673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_12_Left_6674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_12_Left_6675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_12_Left_6676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_12_Left_6677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_12_Left_6678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_12_Left_6679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_12_Left_6680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_12_Left_6681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_12_Left_6682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_12_Left_6683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_12_Left_6684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_12_Left_6685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_12_Left_6686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_12_Left_6687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_12_Left_6688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_12_Left_6689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_12_Left_6690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_12_Left_6691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_12_Left_6692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_12_Left_6693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_12_Left_6694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_12_Left_6695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_12_Left_6696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_12_Left_6697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_12_Left_6698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_12_Left_6699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_12_Left_6700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_12_Left_6701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_12_Left_6702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_12_Left_6703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_12_Left_6704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_12_Left_6705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_12_Left_6706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_12_Left_6707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_12_Left_6708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_12_Left_6709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_12_Left_6710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_12_Left_6711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_12_Left_6712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_12_Left_6713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_12_Left_6714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_12_Left_6715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_12_Left_6716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_12_Left_6717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_12_Left_6718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_12_Left_6719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_12_Left_6720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_12_Left_6721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_12_Left_6722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_12_Left_6723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_12_Left_6724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_12_Left_6725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_12_Left_6726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_12_Left_6727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_12_Left_6728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_12_Left_6729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_12_Left_6730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_12_Left_6731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_12_Left_6732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_12_Left_6733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_12_Left_6734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_12_Left_6735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_12_Left_6736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_12_Left_6737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_12_Left_6738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_12_Left_6739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_12_Left_6740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_12_Left_6741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_12_Left_6742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_12_Left_6743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_12_Left_6744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_12_Left_6745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_12_Left_6746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_12_Left_6747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_12_Left_6748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_12_Left_6749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_12_Left_6750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_12_Left_6751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_12_Left_6752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_12_Left_6753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_12_Left_6754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_12_Left_6755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_12_Left_6756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_12_Left_6757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_12_Left_6758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_12_Left_6759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_12_Left_6760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_12_Left_6761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_12_Left_6762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_12_Left_6763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_12_Left_6764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_12_Left_6765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_12_Left_6766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_12_Left_6767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_12_Left_6768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_12_Left_6769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_12_Left_6770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_12_Left_6771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_12_Left_6772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_12_Left_6773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_12_Left_6774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_12_Left_6775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_12_Left_6776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_12_Left_6777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_12_Left_6778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_12_Left_6779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_12_Left_6780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_12_Left_6781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_12_Left_6782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_12_Left_6783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_12_Left_6784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_12_Left_6785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_12_Left_6786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_12_Left_6787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_12_Left_6788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_12_Left_6789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_12_Left_6790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_12_Left_6791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_12_Left_6792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_12_Left_6793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_12_Left_6794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_12_Left_6795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_12_Left_6796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_12_Left_6797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_12_Left_6798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_12_Left_6799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_12_Left_6800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_12_Left_6801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_12_Left_6802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_12_Left_6803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_12_Right_6804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_12_Right_6805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_12_Right_6806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_12_Right_6807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_12_Right_6808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_12_Right_6809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_12_Right_6810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_12_Right_6811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_12_Right_6812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_12_Right_6813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_12_Right_6814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_12_Right_6815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_12_Right_6816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_12_Right_6817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_12_Right_6818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_12_Right_6819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_12_Right_6820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_12_Right_6821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_12_Right_6822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_12_Right_6823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_12_Right_6824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_12_Right_6825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_12_Right_6826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_12_Right_6827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_12_Right_6828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_12_Right_6829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_12_Right_6830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_12_Right_6831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_12_Right_6832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_12_Right_6833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_12_Right_6834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_12_Right_6835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_12_Right_6836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_12_Right_6837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_12_Right_6838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_12_Right_6839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_12_Right_6840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_12_Right_6841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_12_Right_6842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_12_Right_6843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_12_Right_6844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_12_Right_6845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_12_Right_6846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_12_Right_6847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_12_Right_6848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_12_Right_6849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_12_Right_6850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_12_Right_6851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_12_Right_6852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_12_Right_6853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_12_Right_6854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_12_Right_6855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_12_Right_6856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_12_Right_6857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_12_Right_6858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_12_Right_6859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_12_Right_6860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_12_Right_6861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_12_Right_6862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_12_Right_6863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_12_Right_6864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_12_Right_6865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_12_Right_6866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_12_Right_6867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_12_Right_6868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_12_Right_6869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_12_Right_6870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_12_Right_6871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_12_Right_6872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_12_Right_6873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_12_Right_6874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_12_Right_6875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_12_Right_6876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_12_Right_6877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_12_Right_6878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_12_Right_6879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_12_Right_6880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_12_Right_6881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_12_Right_6882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_12_Right_6883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_12_Right_6884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_12_Right_6885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_12_Right_6886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_12_Right_6887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_12_Right_6888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_12_Right_6889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_12_Right_6890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_12_Right_6891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_12_Right_6892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_12_Right_6893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_12_Right_6894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_12_Right_6895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_12_Right_6896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_12_Right_6897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_12_Right_6898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_12_Right_6899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_12_Right_6900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_12_Right_6901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_12_Right_6902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_12_Right_6903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_12_Right_6904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_12_Right_6905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_12_Right_6906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_12_Right_6907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_12_Right_6908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_12_Right_6909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_12_Right_6910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_12_Right_6911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_12_Right_6912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_12_Right_6913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_12_Right_6914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_12_Right_6915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_12_Right_6916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_12_Right_6917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_12_Right_6918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_12_Right_6919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_12_Right_6920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_12_Right_6921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_12_Right_6922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_12_Right_6923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_12_Right_6924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_12_Right_6925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_12_Right_6926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_12_Right_6927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_12_Right_6928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_12_Right_6929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_12_Right_6930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_12_Right_6931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_12_Right_6932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_12_Right_6933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_12_Right_6934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_12_Right_6935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_12_Right_6936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_12_Right_6937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_12_Right_6938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_12_Right_6939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_12_Right_6940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_12_Right_6941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_12_Right_6942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_12_Right_6943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_12_Right_6944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_12_Right_6945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_12_Right_6946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_12_Right_6947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_12_Right_6948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_12_Right_6949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_12_Right_6950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_12_Right_6951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_12_Right_6952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_12_Right_6953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_12_Right_6954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_12_Right_6955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_12_Right_6956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_12_Right_6957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_12_Right_6958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_12_Right_6959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_12_Right_6960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_12_Right_6961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_12_Right_6962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_12_Right_6963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_12_Right_6964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_12_Right_6965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_12_Right_6966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_12_Right_6967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_12_Right_6968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_12_Right_6969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_12_Right_6970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_12_Right_6971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_12_Right_6972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_12_Right_6973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_12_Right_6974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_12_Right_6975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_12_Right_6976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_12_Right_6977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_12_Right_6978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_12_Right_6979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_12_Right_6980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_12_Right_6981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_12_Right_6982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_12_Right_6983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_12_Right_6984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_12_Right_6985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_12_Right_6986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_12_Right_6987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_12_Right_6988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_12_Right_6989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_12_Right_6990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_12_Right_6991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_12_Right_6992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_12_Right_6993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_12_Right_6994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_12_Right_6995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_12_Right_6996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_12_Right_6997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_12_Right_6998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_12_Right_6999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_12_Right_7000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_12_Right_7001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_12_Right_7002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_12_Right_7003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_12_Right_7004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_12_Right_7005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_12_Right_7006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_12_Right_7007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_12_Right_7008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_12_Right_7009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_12_Right_7010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_12_Right_7011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_12_Right_7012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_12_Right_7013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_12_Right_7014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_12_Right_7015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_12_Right_7016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_12_Right_7017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_12_Right_7018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_12_Right_7019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_12_Right_7020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_12_Right_7021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_12_Right_7022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_12_Right_7023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_12_Right_7024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_12_Right_7025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_12_Right_7026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_12_Right_7027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_12_Right_7028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_12_Right_7029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_12_Right_7030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_12_Right_7031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_12_Right_7032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_12_Right_7033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_12_Right_7034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_12_Right_7035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_12_Right_7036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_12_Right_7037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_12_Right_7038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_12_Right_7039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_12_Right_7040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_12_Right_7041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_12_Right_7042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_12_Right_7043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_12_Right_7044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_12_Right_7045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_12_Right_7046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_12_Right_7047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_12_Right_7048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_12_Right_7049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_12_Right_7050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_12_Right_7051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_12_Right_7052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_12_Right_7053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_12_Right_7054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_12_Right_7055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_12_Right_7056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_12_Right_7057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_12_Right_7058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_12_Right_7059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_12_Right_7060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_12_Right_7061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_12_Right_7062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_12_Right_7063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_12_Right_7064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_12_Right_7065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_12_Right_7066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_12_Right_7067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_12_Right_7068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_12_Right_7069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_12_Right_7070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_12_Right_7071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_12_Right_7072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_12_Right_7073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_12_Right_7074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_12_Right_7075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_12_Right_7076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_12_Right_7077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_12_Right_7078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_12_Right_7079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_12_Right_7080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_12_Right_7081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_12_Right_7082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_12_Right_7083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_12_Right_7084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_12_Right_7085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_12_Right_7086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_12_Right_7087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_12_Right_7088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_12_Right_7089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_12_Right_7090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_12_Right_7091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_12_Right_7092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_12_Right_7093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_12_Right_7094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_12_Right_7095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_12_Right_7096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_12_Right_7097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_12_Right_7098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_12_Right_7099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_12_Right_7100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_12_Right_7101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_12_Right_7102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_12_Right_7103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_12_Right_7104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_12_Right_7105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_12_Right_7106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_12_Right_7107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_12_Right_7108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_12_Right_7109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_12_Right_7110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_12_Right_7111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_12_Right_7112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_12_Right_7113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_12_Right_7114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_12_Right_7115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_12_Right_7116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_12_Right_7117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_12_Right_7118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_12_Right_7119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_12_Right_7120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_12_Right_7121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_12_Right_7122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_12_Right_7123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_12_Right_7124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_12_Right_7125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_12_Right_7126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_12_Right_7127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_13_Left_7128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_13_Left_7129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_13_Left_7130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_13_Left_7131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_13_Left_7132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_13_Left_7133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_13_Left_7134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_13_Left_7135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_13_Left_7136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_13_Left_7137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_13_Left_7138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_13_Left_7139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_13_Left_7140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_13_Left_7141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_13_Left_7142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_13_Left_7143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_13_Left_7144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_13_Left_7145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_13_Left_7146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_13_Left_7147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_13_Left_7148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_13_Left_7149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_13_Left_7150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_13_Left_7151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_13_Left_7152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_13_Left_7153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_13_Left_7154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_13_Left_7155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_13_Left_7156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_13_Left_7157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_13_Left_7158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_13_Left_7159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_13_Left_7160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_13_Left_7161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_13_Left_7162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_13_Left_7163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_13_Left_7164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_13_Left_7165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_13_Left_7166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_13_Left_7167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_13_Left_7168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_13_Left_7169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_13_Left_7170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_13_Left_7171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_13_Left_7172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_13_Left_7173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_13_Left_7174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_13_Left_7175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_13_Left_7176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_13_Left_7177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_13_Left_7178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_13_Left_7179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_13_Left_7180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_13_Left_7181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_13_Left_7182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_13_Left_7183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_13_Left_7184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_13_Left_7185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_13_Left_7186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_13_Left_7187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_13_Left_7188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_13_Left_7189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_13_Left_7190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_13_Left_7191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_13_Left_7192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_13_Left_7193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_13_Left_7194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_13_Left_7195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_13_Left_7196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_13_Left_7197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_13_Left_7198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_13_Left_7199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_13_Left_7200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_13_Left_7201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_13_Left_7202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_13_Left_7203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_13_Left_7204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_13_Left_7205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_13_Left_7206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_13_Left_7207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_13_Left_7208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_13_Left_7209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_13_Left_7210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_13_Left_7211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_13_Left_7212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_13_Left_7213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_13_Left_7214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_13_Left_7215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_13_Left_7216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_13_Left_7217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_13_Left_7218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_13_Left_7219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_13_Left_7220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_13_Left_7221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_13_Left_7222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_13_Left_7223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_13_Left_7224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_13_Left_7225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_13_Left_7226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_13_Left_7227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_13_Left_7228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_13_Left_7229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_13_Left_7230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_13_Left_7231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_13_Left_7232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_13_Left_7233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_13_Left_7234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_13_Left_7235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_13_Left_7236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_13_Left_7237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_13_Left_7238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_13_Left_7239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_13_Left_7240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_13_Left_7241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_13_Left_7242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_13_Left_7243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_13_Left_7244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_13_Left_7245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_13_Left_7246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_13_Left_7247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_13_Left_7248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_13_Left_7249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_13_Left_7250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_13_Left_7251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_13_Left_7252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_13_Left_7253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_13_Left_7254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_13_Left_7255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_13_Left_7256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_13_Left_7257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_13_Left_7258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_13_Left_7259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_13_Left_7260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_13_Left_7261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_13_Left_7262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_13_Left_7263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_13_Left_7264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_13_Left_7265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_13_Left_7266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_13_Left_7267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_13_Left_7268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_13_Left_7269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_13_Left_7270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_13_Left_7271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_13_Left_7272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_13_Left_7273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_13_Left_7274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_13_Left_7275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_13_Left_7276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_13_Left_7277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_13_Left_7278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_13_Left_7279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_13_Left_7280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_13_Left_7281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_13_Left_7282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_13_Left_7283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_13_Left_7284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_13_Left_7285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_13_Left_7286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_13_Left_7287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_13_Left_7288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_13_Left_7289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_13_Left_7290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_13_Left_7291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_13_Left_7292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_13_Left_7293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_13_Left_7294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_13_Left_7295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_13_Left_7296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_13_Left_7297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_13_Left_7298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_13_Left_7299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_13_Left_7300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_13_Left_7301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_13_Left_7302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_13_Left_7303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_13_Left_7304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_13_Left_7305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_13_Left_7306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_13_Left_7307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_13_Left_7308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_13_Left_7309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_13_Left_7310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_13_Left_7311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_13_Left_7312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_13_Left_7313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_13_Left_7314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_13_Left_7315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_13_Left_7316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_13_Left_7317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_13_Left_7318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_13_Left_7319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_13_Left_7320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_13_Left_7321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_13_Left_7322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_13_Left_7323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_13_Left_7324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_13_Left_7325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_13_Left_7326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_13_Left_7327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_13_Left_7328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_13_Left_7329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_13_Left_7330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_13_Left_7331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_13_Left_7332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_13_Left_7333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_13_Left_7334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_13_Left_7335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_13_Left_7336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_13_Left_7337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_13_Left_7338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_13_Left_7339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_13_Left_7340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_13_Left_7341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_13_Left_7342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_13_Left_7343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_13_Left_7344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_13_Left_7345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_13_Left_7346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_13_Left_7347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_13_Left_7348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_13_Left_7349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_13_Left_7350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_13_Left_7351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_13_Left_7352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_13_Left_7353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_13_Left_7354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_13_Left_7355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_13_Left_7356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_13_Left_7357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_13_Left_7358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_13_Left_7359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_13_Left_7360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_13_Left_7361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_13_Left_7362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_13_Left_7363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_13_Left_7364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_13_Left_7365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_13_Left_7366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_13_Left_7367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_13_Left_7368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_13_Left_7369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_13_Left_7370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_13_Left_7371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_13_Left_7372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_13_Left_7373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_13_Left_7374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_13_Left_7375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_13_Left_7376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_13_Left_7377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_13_Left_7378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_13_Left_7379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_13_Left_7380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_13_Left_7381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_13_Left_7382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_13_Left_7383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_13_Left_7384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_13_Left_7385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_13_Left_7386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_13_Left_7387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_13_Left_7388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_13_Left_7389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_13_Left_7390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_13_Left_7391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_13_Left_7392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_13_Left_7393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_13_Left_7394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_13_Left_7395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_13_Left_7396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_13_Left_7397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_13_Left_7398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_13_Left_7399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_13_Left_7400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_13_Left_7401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_13_Left_7402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_13_Left_7403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_13_Left_7404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_13_Left_7405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_13_Left_7406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_13_Left_7407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_13_Left_7408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_13_Left_7409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_13_Left_7410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_13_Left_7411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_13_Left_7412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_13_Left_7413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_13_Left_7414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_13_Left_7415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_13_Left_7416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_13_Left_7417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_13_Left_7418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_13_Left_7419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_13_Left_7420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_13_Left_7421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_13_Left_7422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_13_Left_7423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_13_Left_7424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_13_Left_7425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_13_Left_7426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_13_Left_7427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_13_Left_7428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_13_Left_7429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_13_Left_7430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_13_Left_7431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_13_Left_7432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_13_Left_7433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_13_Left_7434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_13_Left_7435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_13_Left_7436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_13_Left_7437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_13_Left_7438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_13_Left_7439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_13_Left_7440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_13_Left_7441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_13_Left_7442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_13_Left_7443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_13_Left_7444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_13_Left_7445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_13_Left_7446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_13_Left_7447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_13_Left_7448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_13_Left_7449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_13_Left_7450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_13_Left_7451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_13_Right_7452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_13_Right_7453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_13_Right_7454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_13_Right_7455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_13_Right_7456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_13_Right_7457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_13_Right_7458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_13_Right_7459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_13_Right_7460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_13_Right_7461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_13_Right_7462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_13_Right_7463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_13_Right_7464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_13_Right_7465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_13_Right_7466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_13_Right_7467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_13_Right_7468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_13_Right_7469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_13_Right_7470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_13_Right_7471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_13_Right_7472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_13_Right_7473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_13_Right_7474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_13_Right_7475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_13_Right_7476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_13_Right_7477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_13_Right_7478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_13_Right_7479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_13_Right_7480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_13_Right_7481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_13_Right_7482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_13_Right_7483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_13_Right_7484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_13_Right_7485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_13_Right_7486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_13_Right_7487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_13_Right_7488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_13_Right_7489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_13_Right_7490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_13_Right_7491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_13_Right_7492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_13_Right_7493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_13_Right_7494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_13_Right_7495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_13_Right_7496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_13_Right_7497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_13_Right_7498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_13_Right_7499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_13_Right_7500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_13_Right_7501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_13_Right_7502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_13_Right_7503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_13_Right_7504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_13_Right_7505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_13_Right_7506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_13_Right_7507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_13_Right_7508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_13_Right_7509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_13_Right_7510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_13_Right_7511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_13_Right_7512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_13_Right_7513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_13_Right_7514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_13_Right_7515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_13_Right_7516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_13_Right_7517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_13_Right_7518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_13_Right_7519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_13_Right_7520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_13_Right_7521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_13_Right_7522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_13_Right_7523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_13_Right_7524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_13_Right_7525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_13_Right_7526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_13_Right_7527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_13_Right_7528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_13_Right_7529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_13_Right_7530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_13_Right_7531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_13_Right_7532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_13_Right_7533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_13_Right_7534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_13_Right_7535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_13_Right_7536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_13_Right_7537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_13_Right_7538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_13_Right_7539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_13_Right_7540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_13_Right_7541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_13_Right_7542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_13_Right_7543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_13_Right_7544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_13_Right_7545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_13_Right_7546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_13_Right_7547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_13_Right_7548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_13_Right_7549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_13_Right_7550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_13_Right_7551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_13_Right_7552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_13_Right_7553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_13_Right_7554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_13_Right_7555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_13_Right_7556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_13_Right_7557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_13_Right_7558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_13_Right_7559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_13_Right_7560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_13_Right_7561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_13_Right_7562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_13_Right_7563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_13_Right_7564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_13_Right_7565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_13_Right_7566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_13_Right_7567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_13_Right_7568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_13_Right_7569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_13_Right_7570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_13_Right_7571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_13_Right_7572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_13_Right_7573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_13_Right_7574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_13_Right_7575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_13_Right_7576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_13_Right_7577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_13_Right_7578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_13_Right_7579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_13_Right_7580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_13_Right_7581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_13_Right_7582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_13_Right_7583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_13_Right_7584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_13_Right_7585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_13_Right_7586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_13_Right_7587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_13_Right_7588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_13_Right_7589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_13_Right_7590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_13_Right_7591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_13_Right_7592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_13_Right_7593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_13_Right_7594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_13_Right_7595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_13_Right_7596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_13_Right_7597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_13_Right_7598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_13_Right_7599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_13_Right_7600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_13_Right_7601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_13_Right_7602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_13_Right_7603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_13_Right_7604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_13_Right_7605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_13_Right_7606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_13_Right_7607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_13_Right_7608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_13_Right_7609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_13_Right_7610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_13_Right_7611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_13_Right_7612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_13_Right_7613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_13_Right_7614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_13_Right_7615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_13_Right_7616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_13_Right_7617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_13_Right_7618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_13_Right_7619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_13_Right_7620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_13_Right_7621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_13_Right_7622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_13_Right_7623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_13_Right_7624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_13_Right_7625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_13_Right_7626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_13_Right_7627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_13_Right_7628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_13_Right_7629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_13_Right_7630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_13_Right_7631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_13_Right_7632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_13_Right_7633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_13_Right_7634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_13_Right_7635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_13_Right_7636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_13_Right_7637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_13_Right_7638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_13_Right_7639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_13_Right_7640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_13_Right_7641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_13_Right_7642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_13_Right_7643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_13_Right_7644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_13_Right_7645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_13_Right_7646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_13_Right_7647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_13_Right_7648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_13_Right_7649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_13_Right_7650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_13_Right_7651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_13_Right_7652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_13_Right_7653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_13_Right_7654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_13_Right_7655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_13_Right_7656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_13_Right_7657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_13_Right_7658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_13_Right_7659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_13_Right_7660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_13_Right_7661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_13_Right_7662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_13_Right_7663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_13_Right_7664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_13_Right_7665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_13_Right_7666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_13_Right_7667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_13_Right_7668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_13_Right_7669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_13_Right_7670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_13_Right_7671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_13_Right_7672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_13_Right_7673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_13_Right_7674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_13_Right_7675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_13_Right_7676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_13_Right_7677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_13_Right_7678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_13_Right_7679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_13_Right_7680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_13_Right_7681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_13_Right_7682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_13_Right_7683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_13_Right_7684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_13_Right_7685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_13_Right_7686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_13_Right_7687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_13_Right_7688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_13_Right_7689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_13_Right_7690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_13_Right_7691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_13_Right_7692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_13_Right_7693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_13_Right_7694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_13_Right_7695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_13_Right_7696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_13_Right_7697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_13_Right_7698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_13_Right_7699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_13_Right_7700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_13_Right_7701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_13_Right_7702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_13_Right_7703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_13_Right_7704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_13_Right_7705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_13_Right_7706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_13_Right_7707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_13_Right_7708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_13_Right_7709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_13_Right_7710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_13_Right_7711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_13_Right_7712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_13_Right_7713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_13_Right_7714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_13_Right_7715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_13_Right_7716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_13_Right_7717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_13_Right_7718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_13_Right_7719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_13_Right_7720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_13_Right_7721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_13_Right_7722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_13_Right_7723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_13_Right_7724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_13_Right_7725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_13_Right_7726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_13_Right_7727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_13_Right_7728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_13_Right_7729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_13_Right_7730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_13_Right_7731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_13_Right_7732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_13_Right_7733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_13_Right_7734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_13_Right_7735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_13_Right_7736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_13_Right_7737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_13_Right_7738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_13_Right_7739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_13_Right_7740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_13_Right_7741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_13_Right_7742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_13_Right_7743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_13_Right_7744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_13_Right_7745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_13_Right_7746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_13_Right_7747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_13_Right_7748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_13_Right_7749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_13_Right_7750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_13_Right_7751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_13_Right_7752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_13_Right_7753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_13_Right_7754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_13_Right_7755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_13_Right_7756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_13_Right_7757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_13_Right_7758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_13_Right_7759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_13_Right_7760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_13_Right_7761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_13_Right_7762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_13_Right_7763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_13_Right_7764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_13_Right_7765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_13_Right_7766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_13_Right_7767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_13_Right_7768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_13_Right_7769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_13_Right_7770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_13_Right_7771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_13_Right_7772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_13_Right_7773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_13_Right_7774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_13_Right_7775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_14_Left_7776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_14_Left_7777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_14_Left_7778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_14_Left_7779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_14_Left_7780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_14_Left_7781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_14_Left_7782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_14_Left_7783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_14_Left_7784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_14_Left_7785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_14_Left_7786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_14_Left_7787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_14_Left_7788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_14_Left_7789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_14_Left_7790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_14_Left_7791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_14_Left_7792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_14_Left_7793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_14_Left_7794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_14_Left_7795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_14_Left_7796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_14_Left_7797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_14_Left_7798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_14_Left_7799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_14_Left_7800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_14_Left_7801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_14_Left_7802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_14_Left_7803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_14_Left_7804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_14_Left_7805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_14_Left_7806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_14_Left_7807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_14_Left_7808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_14_Left_7809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_14_Left_7810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_14_Left_7811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_14_Left_7812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_14_Left_7813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_14_Left_7814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_14_Left_7815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_14_Left_7816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_14_Left_7817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_14_Left_7818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_14_Left_7819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_14_Left_7820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_14_Left_7821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_14_Left_7822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_14_Left_7823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_14_Left_7824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_14_Left_7825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_14_Left_7826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_14_Left_7827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_14_Left_7828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_14_Left_7829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_14_Left_7830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_14_Left_7831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_14_Left_7832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_14_Left_7833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_14_Left_7834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_14_Left_7835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_14_Left_7836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_14_Left_7837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_14_Left_7838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_14_Left_7839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_14_Left_7840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_14_Left_7841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_14_Left_7842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_14_Left_7843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_14_Left_7844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_14_Left_7845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_14_Left_7846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_14_Left_7847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_14_Left_7848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_14_Left_7849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_14_Left_7850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_14_Left_7851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_14_Left_7852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_14_Left_7853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_14_Left_7854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_14_Left_7855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_14_Left_7856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_14_Left_7857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_14_Left_7858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_14_Left_7859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_14_Left_7860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_14_Left_7861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_14_Left_7862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_14_Left_7863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_14_Left_7864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_14_Left_7865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_14_Left_7866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_14_Left_7867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_14_Left_7868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_14_Left_7869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_14_Left_7870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_14_Left_7871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_14_Left_7872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_14_Left_7873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_14_Left_7874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_14_Left_7875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_14_Left_7876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_14_Left_7877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_14_Left_7878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_14_Left_7879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_14_Left_7880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_14_Left_7881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_14_Left_7882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_14_Left_7883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_14_Left_7884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_14_Left_7885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_14_Left_7886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_14_Left_7887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_14_Left_7888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_14_Left_7889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_14_Left_7890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_14_Left_7891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_14_Left_7892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_14_Left_7893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_14_Left_7894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_14_Left_7895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_14_Left_7896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_14_Left_7897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_14_Left_7898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_14_Left_7899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_14_Left_7900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_14_Left_7901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_14_Left_7902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_14_Left_7903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_14_Left_7904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_14_Left_7905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_14_Left_7906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_14_Left_7907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_14_Left_7908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_14_Left_7909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_14_Left_7910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_14_Left_7911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_14_Left_7912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_14_Left_7913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_14_Left_7914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_14_Left_7915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_14_Left_7916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_14_Left_7917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_14_Left_7918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_14_Left_7919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_14_Left_7920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_14_Left_7921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_14_Left_7922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_14_Left_7923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_14_Left_7924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_14_Left_7925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_14_Left_7926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_14_Left_7927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_14_Left_7928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_14_Left_7929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_14_Left_7930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_14_Left_7931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_14_Left_7932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_14_Left_7933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_14_Left_7934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_14_Left_7935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_14_Left_7936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_14_Left_7937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_14_Left_7938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_14_Left_7939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_14_Left_7940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_14_Left_7941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_14_Left_7942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_14_Left_7943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_14_Left_7944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_14_Left_7945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_14_Left_7946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_14_Left_7947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_14_Left_7948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_14_Left_7949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_14_Left_7950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_14_Left_7951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_14_Left_7952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_14_Left_7953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_14_Left_7954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_14_Left_7955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_14_Left_7956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_14_Left_7957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_14_Left_7958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_14_Left_7959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_14_Left_7960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_14_Left_7961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_14_Left_7962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_14_Left_7963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_14_Left_7964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_14_Left_7965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_14_Left_7966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_14_Left_7967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_14_Left_7968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_14_Left_7969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_14_Left_7970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_14_Left_7971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_14_Left_7972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_14_Left_7973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_14_Left_7974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_14_Left_7975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_14_Left_7976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_14_Left_7977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_14_Left_7978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_14_Left_7979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_14_Left_7980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_14_Left_7981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_14_Left_7982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_14_Left_7983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_14_Left_7984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_14_Left_7985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_14_Left_7986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_14_Left_7987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_14_Left_7988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_14_Left_7989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_14_Left_7990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_14_Left_7991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_14_Left_7992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_14_Left_7993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_14_Left_7994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_14_Left_7995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_14_Left_7996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_14_Left_7997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_14_Left_7998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_14_Left_7999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_14_Left_8000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_14_Left_8001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_14_Left_8002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_14_Left_8003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_14_Left_8004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_14_Left_8005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_14_Left_8006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_14_Left_8007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_14_Left_8008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_14_Left_8009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_14_Left_8010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_14_Left_8011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_14_Left_8012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_14_Left_8013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_14_Left_8014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_14_Left_8015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_14_Left_8016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_14_Left_8017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_14_Left_8018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_14_Left_8019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_14_Left_8020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_14_Left_8021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_14_Left_8022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_14_Left_8023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_14_Left_8024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_14_Left_8025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_14_Left_8026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_14_Left_8027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_14_Left_8028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_14_Left_8029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_14_Left_8030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_14_Left_8031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_14_Left_8032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_14_Left_8033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_14_Left_8034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_14_Left_8035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_14_Left_8036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_14_Left_8037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_14_Left_8038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_14_Left_8039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_14_Left_8040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_14_Left_8041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_14_Left_8042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_14_Left_8043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_14_Left_8044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_14_Left_8045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_14_Left_8046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_14_Left_8047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_14_Left_8048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_14_Left_8049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_14_Left_8050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_14_Left_8051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_14_Left_8052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_14_Left_8053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_14_Left_8054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_14_Left_8055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_14_Left_8056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_14_Left_8057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_14_Left_8058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_14_Left_8059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_14_Left_8060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_14_Left_8061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_14_Left_8062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_14_Left_8063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_14_Left_8064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_14_Left_8065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_14_Left_8066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_14_Left_8067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_14_Left_8068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_14_Left_8069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_14_Left_8070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_14_Left_8071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_14_Left_8072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_14_Left_8073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_14_Left_8074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_14_Left_8075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_14_Left_8076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_14_Left_8077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_14_Left_8078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_14_Left_8079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_14_Left_8080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_14_Left_8081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_14_Left_8082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_14_Left_8083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_14_Left_8084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_14_Left_8085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_14_Left_8086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_14_Left_8087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_14_Left_8088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_14_Left_8089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_14_Left_8090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_14_Left_8091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_14_Left_8092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_14_Left_8093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_14_Left_8094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_14_Left_8095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_14_Left_8096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_14_Left_8097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_14_Left_8098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_14_Left_8099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_14_Right_8100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_14_Right_8101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_14_Right_8102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_14_Right_8103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_14_Right_8104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_14_Right_8105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_14_Right_8106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_14_Right_8107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_14_Right_8108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_14_Right_8109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_14_Right_8110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_14_Right_8111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_14_Right_8112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_14_Right_8113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_14_Right_8114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_14_Right_8115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_14_Right_8116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_14_Right_8117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_14_Right_8118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_14_Right_8119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_14_Right_8120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_14_Right_8121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_14_Right_8122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_14_Right_8123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_14_Right_8124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_14_Right_8125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_14_Right_8126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_14_Right_8127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_14_Right_8128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_14_Right_8129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_14_Right_8130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_14_Right_8131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_14_Right_8132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_14_Right_8133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_14_Right_8134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_14_Right_8135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_14_Right_8136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_14_Right_8137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_14_Right_8138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_14_Right_8139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_14_Right_8140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_14_Right_8141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_14_Right_8142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_14_Right_8143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_14_Right_8144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_14_Right_8145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_14_Right_8146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_14_Right_8147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_14_Right_8148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_14_Right_8149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_14_Right_8150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_14_Right_8151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_14_Right_8152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_14_Right_8153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_14_Right_8154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_14_Right_8155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_14_Right_8156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_14_Right_8157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_14_Right_8158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_14_Right_8159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_14_Right_8160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_14_Right_8161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_14_Right_8162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_14_Right_8163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_14_Right_8164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_14_Right_8165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_14_Right_8166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_14_Right_8167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_14_Right_8168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_14_Right_8169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_14_Right_8170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_14_Right_8171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_14_Right_8172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_14_Right_8173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_14_Right_8174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_14_Right_8175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_14_Right_8176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_14_Right_8177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_14_Right_8178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_14_Right_8179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_14_Right_8180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_14_Right_8181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_14_Right_8182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_14_Right_8183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_14_Right_8184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_14_Right_8185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_14_Right_8186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_14_Right_8187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_14_Right_8188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_14_Right_8189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_14_Right_8190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_14_Right_8191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_14_Right_8192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_14_Right_8193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_14_Right_8194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_14_Right_8195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_14_Right_8196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_14_Right_8197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_14_Right_8198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_14_Right_8199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_14_Right_8200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_14_Right_8201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_14_Right_8202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_14_Right_8203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_14_Right_8204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_14_Right_8205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_14_Right_8206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_14_Right_8207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_14_Right_8208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_14_Right_8209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_14_Right_8210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_14_Right_8211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_14_Right_8212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_14_Right_8213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_14_Right_8214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_14_Right_8215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_14_Right_8216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_14_Right_8217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_14_Right_8218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_14_Right_8219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_14_Right_8220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_14_Right_8221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_14_Right_8222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_14_Right_8223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_14_Right_8224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_14_Right_8225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_14_Right_8226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_14_Right_8227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_14_Right_8228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_14_Right_8229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_14_Right_8230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_14_Right_8231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_14_Right_8232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_14_Right_8233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_14_Right_8234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_14_Right_8235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_14_Right_8236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_14_Right_8237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_14_Right_8238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_14_Right_8239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_14_Right_8240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_14_Right_8241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_14_Right_8242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_14_Right_8243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_14_Right_8244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_14_Right_8245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_14_Right_8246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_14_Right_8247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_14_Right_8248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_14_Right_8249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_14_Right_8250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_14_Right_8251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_14_Right_8252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_14_Right_8253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_14_Right_8254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_14_Right_8255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_14_Right_8256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_14_Right_8257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_14_Right_8258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_14_Right_8259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_14_Right_8260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_14_Right_8261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_14_Right_8262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_14_Right_8263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_14_Right_8264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_14_Right_8265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_14_Right_8266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_14_Right_8267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_14_Right_8268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_14_Right_8269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_14_Right_8270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_14_Right_8271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_14_Right_8272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_14_Right_8273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_14_Right_8274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_14_Right_8275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_14_Right_8276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_14_Right_8277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_14_Right_8278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_14_Right_8279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_14_Right_8280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_14_Right_8281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_14_Right_8282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_14_Right_8283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_14_Right_8284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_14_Right_8285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_14_Right_8286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_14_Right_8287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_14_Right_8288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_14_Right_8289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_14_Right_8290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_14_Right_8291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_14_Right_8292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_14_Right_8293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_14_Right_8294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_14_Right_8295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_14_Right_8296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_14_Right_8297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_14_Right_8298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_14_Right_8299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_14_Right_8300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_14_Right_8301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_14_Right_8302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_14_Right_8303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_14_Right_8304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_14_Right_8305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_14_Right_8306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_14_Right_8307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_14_Right_8308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_14_Right_8309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_14_Right_8310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_14_Right_8311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_14_Right_8312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_14_Right_8313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_14_Right_8314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_14_Right_8315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_14_Right_8316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_14_Right_8317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_14_Right_8318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_14_Right_8319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_14_Right_8320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_14_Right_8321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_14_Right_8322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_14_Right_8323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_14_Right_8324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_14_Right_8325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_14_Right_8326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_14_Right_8327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_14_Right_8328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_14_Right_8329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_14_Right_8330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_14_Right_8331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_14_Right_8332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_14_Right_8333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_14_Right_8334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_14_Right_8335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_14_Right_8336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_14_Right_8337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_14_Right_8338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_14_Right_8339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_14_Right_8340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_14_Right_8341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_14_Right_8342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_14_Right_8343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_14_Right_8344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_14_Right_8345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_14_Right_8346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_14_Right_8347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_14_Right_8348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_14_Right_8349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_14_Right_8350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_14_Right_8351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_14_Right_8352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_14_Right_8353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_14_Right_8354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_14_Right_8355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_14_Right_8356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_14_Right_8357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_14_Right_8358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_14_Right_8359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_14_Right_8360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_14_Right_8361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_14_Right_8362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_14_Right_8363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_14_Right_8364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_14_Right_8365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_14_Right_8366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_14_Right_8367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_14_Right_8368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_14_Right_8369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_14_Right_8370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_14_Right_8371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_14_Right_8372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_14_Right_8373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_14_Right_8374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_14_Right_8375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_14_Right_8376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_14_Right_8377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_14_Right_8378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_14_Right_8379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_14_Right_8380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_14_Right_8381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_14_Right_8382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_14_Right_8383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_14_Right_8384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_14_Right_8385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_14_Right_8386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_14_Right_8387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_14_Right_8388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_14_Right_8389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_14_Right_8390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_14_Right_8391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_14_Right_8392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_14_Right_8393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_14_Right_8394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_14_Right_8395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_14_Right_8396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_14_Right_8397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_14_Right_8398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_14_Right_8399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_14_Right_8400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_14_Right_8401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_14_Right_8402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_14_Right_8403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_14_Right_8404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_14_Right_8405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_14_Right_8406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_14_Right_8407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_14_Right_8408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_14_Right_8409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_14_Right_8410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_14_Right_8411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_14_Right_8412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_14_Right_8413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_14_Right_8414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_14_Right_8415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_14_Right_8416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_14_Right_8417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_14_Right_8418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_14_Right_8419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_14_Right_8420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_14_Right_8421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_14_Right_8422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_14_Right_8423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_15_Left_8424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_15_Left_8425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_15_Left_8426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_15_Left_8427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_15_Left_8428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_15_Left_8429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_15_Left_8430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_15_Left_8431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_15_Left_8432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_15_Left_8433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_15_Left_8434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_15_Left_8435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_15_Left_8436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_15_Left_8437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_15_Left_8438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_15_Left_8439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_15_Left_8440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_15_Left_8441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_15_Left_8442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_15_Left_8443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_15_Left_8444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_15_Left_8445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_15_Left_8446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_15_Left_8447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_15_Left_8448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_15_Left_8449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_15_Left_8450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_15_Left_8451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_15_Left_8452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_15_Left_8453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_15_Left_8454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_15_Left_8455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_15_Left_8456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_15_Left_8457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_15_Left_8458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_15_Left_8459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_15_Left_8460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_15_Left_8461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_15_Left_8462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_15_Left_8463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_15_Left_8464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_15_Left_8465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_15_Left_8466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_15_Left_8467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_15_Left_8468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_15_Left_8469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_15_Left_8470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_15_Left_8471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_15_Left_8472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_15_Left_8473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_15_Left_8474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_15_Left_8475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_15_Left_8476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_15_Left_8477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_15_Left_8478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_15_Left_8479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_15_Left_8480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_15_Left_8481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_15_Left_8482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_15_Left_8483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_15_Left_8484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_15_Left_8485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_15_Left_8486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_15_Left_8487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_15_Left_8488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_15_Left_8489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_15_Left_8490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_15_Left_8491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_15_Left_8492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_15_Left_8493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_15_Left_8494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_15_Left_8495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_15_Left_8496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_15_Left_8497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_15_Left_8498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_15_Left_8499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_15_Left_8500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_15_Left_8501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_15_Left_8502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_15_Left_8503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_15_Left_8504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_15_Left_8505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_15_Left_8506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_15_Left_8507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_15_Left_8508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_15_Left_8509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_15_Left_8510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_15_Left_8511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_15_Left_8512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_15_Left_8513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_15_Left_8514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_15_Left_8515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_15_Left_8516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_15_Left_8517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_15_Left_8518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_15_Left_8519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_15_Left_8520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_15_Left_8521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_15_Left_8522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_15_Left_8523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_15_Left_8524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_15_Left_8525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_15_Left_8526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_15_Left_8527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_15_Left_8528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_15_Left_8529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_15_Left_8530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_15_Left_8531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_15_Left_8532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_15_Left_8533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_15_Left_8534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_15_Left_8535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_15_Left_8536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_15_Left_8537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_15_Left_8538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_15_Left_8539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_15_Left_8540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_15_Left_8541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_15_Left_8542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_15_Left_8543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_15_Left_8544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_15_Left_8545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_15_Left_8546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_15_Left_8547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_15_Left_8548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_15_Left_8549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_15_Left_8550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_15_Left_8551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_15_Left_8552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_15_Left_8553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_15_Left_8554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_15_Left_8555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_15_Left_8556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_15_Left_8557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_15_Left_8558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_15_Left_8559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_15_Left_8560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_15_Left_8561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_15_Left_8562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_15_Left_8563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_15_Left_8564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_15_Left_8565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_15_Left_8566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_15_Left_8567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_15_Left_8568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_15_Left_8569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_15_Left_8570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_15_Left_8571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_15_Left_8572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_15_Left_8573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_15_Left_8574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_15_Left_8575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_15_Left_8576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_15_Left_8577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_15_Left_8578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_15_Left_8579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_15_Left_8580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_15_Left_8581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_15_Left_8582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_15_Left_8583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_15_Left_8584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_15_Left_8585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_15_Left_8586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_15_Left_8587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_15_Left_8588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_15_Left_8589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_15_Left_8590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_15_Left_8591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_15_Left_8592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_15_Left_8593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_15_Left_8594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_15_Left_8595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_15_Left_8596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_15_Left_8597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_15_Left_8598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_15_Left_8599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_15_Left_8600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_15_Left_8601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_15_Left_8602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_15_Left_8603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_15_Left_8604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_15_Left_8605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_15_Left_8606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_15_Left_8607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_15_Left_8608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_15_Left_8609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_15_Left_8610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_15_Left_8611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_15_Left_8612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_15_Left_8613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_15_Left_8614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_15_Left_8615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_15_Left_8616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_15_Left_8617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_15_Left_8618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_15_Left_8619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_15_Left_8620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_15_Left_8621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_15_Left_8622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_15_Left_8623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_15_Left_8624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_15_Left_8625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_15_Left_8626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_15_Left_8627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_15_Left_8628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_15_Left_8629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_15_Left_8630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_15_Left_8631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_15_Left_8632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_15_Left_8633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_15_Left_8634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_15_Left_8635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_15_Left_8636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_15_Left_8637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_15_Left_8638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_15_Left_8639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_15_Left_8640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_15_Left_8641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_15_Left_8642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_15_Left_8643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_15_Left_8644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_15_Left_8645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_15_Left_8646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_15_Left_8647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_15_Left_8648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_15_Left_8649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_15_Left_8650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_15_Left_8651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_15_Left_8652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_15_Left_8653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_15_Left_8654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_15_Left_8655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_15_Left_8656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_15_Left_8657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_15_Left_8658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_15_Left_8659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_15_Left_8660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_15_Left_8661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_15_Left_8662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_15_Left_8663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_15_Left_8664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_15_Left_8665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_15_Left_8666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_15_Left_8667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_15_Left_8668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_15_Left_8669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_15_Left_8670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_15_Left_8671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_15_Left_8672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_15_Left_8673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_15_Left_8674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_15_Left_8675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_15_Left_8676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_15_Left_8677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_15_Left_8678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_15_Left_8679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_15_Left_8680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_15_Left_8681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_15_Left_8682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_15_Left_8683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_15_Left_8684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_15_Left_8685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_15_Left_8686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_15_Left_8687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_15_Left_8688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_15_Left_8689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_15_Left_8690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_15_Left_8691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_15_Left_8692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_15_Left_8693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_15_Left_8694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_15_Left_8695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_15_Left_8696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_15_Left_8697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_15_Left_8698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_15_Left_8699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_15_Left_8700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_15_Left_8701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_15_Left_8702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_15_Left_8703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_15_Left_8704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_15_Left_8705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_15_Left_8706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_15_Left_8707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_15_Left_8708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_15_Left_8709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_15_Left_8710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_15_Left_8711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_15_Left_8712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_15_Left_8713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_15_Left_8714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_15_Left_8715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_15_Left_8716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_15_Left_8717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_15_Left_8718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_15_Left_8719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_15_Left_8720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_15_Left_8721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_15_Left_8722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_15_Left_8723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_15_Left_8724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_15_Left_8725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_15_Left_8726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_15_Left_8727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_15_Left_8728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_15_Left_8729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_15_Left_8730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_15_Left_8731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_15_Left_8732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_15_Left_8733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_15_Left_8734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_15_Left_8735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_15_Left_8736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_15_Left_8737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_15_Left_8738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_15_Left_8739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_15_Left_8740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_15_Left_8741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_15_Left_8742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_15_Left_8743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_15_Left_8744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_15_Left_8745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_15_Left_8746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_15_Left_8747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_15_Right_8748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_15_Right_8749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_15_Right_8750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_15_Right_8751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_15_Right_8752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_15_Right_8753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_15_Right_8754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_15_Right_8755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_15_Right_8756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_15_Right_8757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_15_Right_8758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_15_Right_8759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_15_Right_8760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_15_Right_8761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_15_Right_8762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_15_Right_8763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_15_Right_8764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_15_Right_8765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_15_Right_8766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_15_Right_8767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_15_Right_8768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_15_Right_8769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_15_Right_8770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_15_Right_8771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_15_Right_8772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_15_Right_8773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_15_Right_8774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_15_Right_8775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_15_Right_8776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_15_Right_8777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_15_Right_8778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_15_Right_8779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_15_Right_8780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_15_Right_8781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_15_Right_8782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_15_Right_8783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_15_Right_8784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_15_Right_8785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_15_Right_8786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_15_Right_8787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_15_Right_8788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_15_Right_8789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_15_Right_8790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_15_Right_8791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_15_Right_8792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_15_Right_8793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_15_Right_8794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_15_Right_8795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_15_Right_8796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_15_Right_8797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_15_Right_8798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_15_Right_8799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_15_Right_8800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_15_Right_8801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_15_Right_8802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_15_Right_8803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_15_Right_8804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_15_Right_8805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_15_Right_8806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_15_Right_8807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_15_Right_8808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_15_Right_8809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_15_Right_8810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_15_Right_8811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_15_Right_8812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_15_Right_8813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_15_Right_8814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_15_Right_8815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_15_Right_8816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_15_Right_8817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_15_Right_8818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_15_Right_8819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_15_Right_8820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_15_Right_8821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_15_Right_8822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_15_Right_8823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_15_Right_8824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_15_Right_8825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_15_Right_8826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_15_Right_8827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_15_Right_8828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_15_Right_8829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_15_Right_8830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_15_Right_8831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_15_Right_8832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_15_Right_8833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_15_Right_8834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_15_Right_8835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_15_Right_8836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_15_Right_8837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_15_Right_8838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_15_Right_8839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_15_Right_8840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_15_Right_8841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_15_Right_8842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_15_Right_8843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_15_Right_8844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_15_Right_8845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_15_Right_8846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_15_Right_8847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_15_Right_8848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_15_Right_8849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_15_Right_8850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_15_Right_8851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_15_Right_8852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_15_Right_8853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_15_Right_8854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_15_Right_8855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_15_Right_8856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_15_Right_8857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_15_Right_8858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_15_Right_8859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_15_Right_8860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_15_Right_8861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_15_Right_8862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_15_Right_8863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_15_Right_8864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_15_Right_8865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_15_Right_8866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_15_Right_8867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_15_Right_8868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_15_Right_8869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_15_Right_8870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_15_Right_8871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_15_Right_8872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_15_Right_8873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_15_Right_8874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_15_Right_8875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_15_Right_8876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_15_Right_8877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_15_Right_8878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_15_Right_8879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_15_Right_8880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_15_Right_8881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_15_Right_8882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_15_Right_8883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_15_Right_8884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_15_Right_8885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_15_Right_8886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_15_Right_8887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_15_Right_8888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_15_Right_8889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_15_Right_8890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_15_Right_8891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_15_Right_8892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_15_Right_8893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_15_Right_8894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_15_Right_8895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_15_Right_8896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_15_Right_8897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_15_Right_8898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_15_Right_8899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_15_Right_8900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_15_Right_8901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_15_Right_8902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_15_Right_8903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_15_Right_8904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_15_Right_8905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_15_Right_8906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_15_Right_8907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_15_Right_8908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_15_Right_8909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_15_Right_8910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_15_Right_8911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_15_Right_8912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_15_Right_8913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_15_Right_8914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_15_Right_8915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_15_Right_8916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_15_Right_8917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_15_Right_8918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_15_Right_8919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_15_Right_8920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_15_Right_8921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_15_Right_8922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_15_Right_8923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_15_Right_8924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_15_Right_8925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_15_Right_8926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_15_Right_8927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_15_Right_8928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_15_Right_8929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_15_Right_8930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_15_Right_8931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_15_Right_8932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_15_Right_8933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_15_Right_8934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_15_Right_8935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_15_Right_8936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_15_Right_8937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_15_Right_8938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_15_Right_8939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_15_Right_8940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_15_Right_8941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_15_Right_8942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_15_Right_8943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_15_Right_8944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_15_Right_8945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_15_Right_8946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_15_Right_8947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_15_Right_8948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_15_Right_8949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_15_Right_8950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_15_Right_8951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_15_Right_8952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_15_Right_8953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_15_Right_8954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_15_Right_8955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_15_Right_8956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_15_Right_8957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_15_Right_8958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_15_Right_8959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_15_Right_8960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_15_Right_8961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_15_Right_8962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_15_Right_8963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_15_Right_8964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_15_Right_8965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_15_Right_8966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_15_Right_8967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_15_Right_8968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_15_Right_8969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_15_Right_8970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_15_Right_8971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_15_Right_8972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_15_Right_8973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_15_Right_8974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_15_Right_8975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_15_Right_8976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_15_Right_8977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_15_Right_8978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_15_Right_8979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_15_Right_8980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_15_Right_8981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_15_Right_8982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_15_Right_8983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_15_Right_8984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_15_Right_8985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_15_Right_8986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_15_Right_8987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_15_Right_8988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_15_Right_8989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_15_Right_8990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_15_Right_8991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_15_Right_8992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_15_Right_8993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_15_Right_8994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_15_Right_8995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_15_Right_8996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_15_Right_8997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_15_Right_8998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_15_Right_8999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_15_Right_9000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_15_Right_9001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_15_Right_9002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_15_Right_9003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_15_Right_9004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_15_Right_9005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_15_Right_9006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_15_Right_9007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_15_Right_9008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_15_Right_9009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_15_Right_9010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_15_Right_9011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_15_Right_9012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_15_Right_9013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_15_Right_9014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_15_Right_9015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_15_Right_9016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_15_Right_9017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_15_Right_9018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_15_Right_9019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_15_Right_9020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_15_Right_9021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_15_Right_9022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_15_Right_9023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_15_Right_9024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_15_Right_9025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_15_Right_9026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_15_Right_9027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_15_Right_9028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_15_Right_9029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_15_Right_9030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_15_Right_9031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_15_Right_9032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_15_Right_9033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_15_Right_9034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_15_Right_9035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_15_Right_9036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_15_Right_9037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_15_Right_9038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_15_Right_9039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_15_Right_9040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_15_Right_9041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_15_Right_9042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_15_Right_9043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_15_Right_9044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_15_Right_9045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_15_Right_9046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_15_Right_9047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_15_Right_9048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_15_Right_9049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_15_Right_9050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_15_Right_9051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_15_Right_9052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_15_Right_9053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_15_Right_9054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_15_Right_9055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_15_Right_9056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_15_Right_9057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_15_Right_9058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_15_Right_9059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_15_Right_9060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_15_Right_9061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_15_Right_9062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_15_Right_9063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_15_Right_9064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_15_Right_9065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_15_Right_9066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_15_Right_9067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_15_Right_9068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_15_Right_9069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_15_Right_9070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_15_Right_9071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_16_Left_9072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_16_Left_9073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_16_Left_9074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_16_Left_9075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_16_Left_9076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_16_Left_9077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_16_Left_9078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_16_Left_9079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_16_Left_9080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_16_Left_9081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_16_Left_9082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_16_Left_9083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_16_Left_9084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_16_Left_9085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_16_Left_9086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_16_Left_9087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_16_Left_9088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_16_Left_9089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_16_Left_9090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_16_Left_9091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_16_Left_9092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_16_Left_9093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_16_Left_9094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_16_Left_9095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_16_Left_9096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_16_Left_9097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_16_Left_9098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_16_Left_9099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_16_Left_9100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_16_Left_9101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_16_Left_9102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_16_Left_9103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_16_Left_9104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_16_Left_9105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_16_Left_9106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_16_Left_9107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_16_Left_9108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_16_Left_9109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_16_Left_9110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_16_Left_9111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_16_Left_9112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_16_Left_9113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_16_Left_9114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_16_Left_9115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_16_Left_9116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_16_Left_9117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_16_Left_9118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_16_Left_9119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_16_Left_9120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_16_Left_9121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_16_Left_9122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_16_Left_9123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_16_Left_9124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_16_Left_9125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_16_Left_9126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_16_Left_9127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_16_Left_9128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_16_Left_9129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_16_Left_9130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_16_Left_9131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_16_Left_9132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_16_Left_9133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_16_Left_9134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_16_Left_9135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_16_Left_9136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_16_Left_9137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_16_Left_9138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_16_Left_9139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_16_Left_9140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_16_Left_9141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_16_Left_9142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_16_Left_9143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_16_Left_9144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_16_Left_9145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_16_Left_9146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_16_Left_9147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_16_Left_9148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_16_Left_9149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_16_Left_9150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_16_Left_9151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_16_Left_9152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_16_Left_9153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_16_Left_9154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_16_Left_9155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_16_Left_9156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_16_Left_9157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_16_Left_9158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_16_Left_9159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_16_Left_9160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_16_Left_9161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_16_Left_9162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_16_Left_9163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_16_Left_9164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_16_Left_9165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_16_Left_9166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_16_Left_9167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_16_Left_9168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_16_Left_9169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_16_Left_9170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_16_Left_9171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_16_Left_9172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_16_Left_9173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_16_Left_9174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_16_Left_9175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_16_Left_9176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_16_Left_9177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_16_Left_9178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_16_Left_9179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_16_Left_9180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_16_Left_9181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_16_Left_9182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_16_Left_9183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_16_Left_9184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_16_Left_9185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_16_Left_9186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_16_Left_9187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_16_Left_9188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_16_Left_9189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_16_Left_9190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_16_Left_9191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_16_Left_9192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_16_Left_9193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_16_Left_9194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_16_Left_9195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_16_Left_9196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_16_Left_9197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_16_Left_9198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_16_Left_9199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_16_Left_9200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_16_Left_9201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_16_Left_9202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_16_Left_9203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_16_Left_9204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_16_Left_9205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_16_Left_9206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_16_Left_9207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_16_Left_9208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_16_Left_9209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_16_Left_9210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_16_Left_9211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_16_Left_9212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_16_Left_9213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_16_Left_9214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_16_Left_9215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_16_Left_9216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_16_Left_9217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_16_Left_9218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_16_Left_9219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_16_Left_9220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_16_Left_9221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_16_Left_9222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_16_Left_9223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_16_Left_9224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_16_Left_9225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_16_Left_9226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_16_Left_9227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_16_Left_9228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_16_Left_9229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_16_Left_9230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_16_Left_9231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_16_Left_9232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_16_Left_9233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_16_Left_9234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_16_Left_9235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_16_Left_9236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_16_Left_9237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_16_Left_9238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_16_Left_9239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_16_Left_9240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_16_Left_9241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_16_Left_9242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_16_Left_9243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_16_Left_9244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_16_Left_9245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_16_Left_9246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_16_Left_9247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_16_Left_9248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_16_Left_9249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_16_Left_9250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_16_Left_9251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_16_Left_9252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_16_Left_9253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_16_Left_9254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_16_Left_9255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_16_Left_9256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_16_Left_9257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_16_Left_9258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_16_Left_9259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_16_Left_9260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_16_Left_9261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_16_Left_9262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_16_Left_9263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_16_Left_9264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_16_Left_9265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_16_Left_9266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_16_Left_9267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_16_Left_9268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_16_Left_9269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_16_Left_9270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_16_Left_9271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_16_Left_9272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_16_Left_9273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_16_Left_9274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_16_Left_9275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_16_Left_9276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_16_Left_9277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_16_Left_9278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_16_Left_9279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_16_Left_9280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_16_Left_9281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_16_Left_9282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_16_Left_9283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_16_Left_9284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_16_Left_9285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_16_Left_9286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_16_Left_9287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_16_Left_9288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_16_Left_9289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_16_Left_9290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_16_Left_9291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_16_Left_9292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_16_Left_9293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_16_Left_9294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_16_Left_9295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_16_Left_9296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_16_Left_9297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_16_Left_9298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_16_Left_9299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_16_Left_9300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_16_Left_9301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_16_Left_9302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_16_Left_9303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_16_Left_9304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_16_Left_9305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_16_Left_9306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_16_Left_9307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_16_Left_9308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_16_Left_9309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_16_Left_9310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_16_Left_9311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_16_Left_9312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_16_Left_9313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_16_Left_9314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_16_Left_9315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_16_Left_9316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_16_Left_9317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_16_Left_9318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_16_Left_9319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_16_Left_9320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_16_Left_9321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_16_Left_9322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_16_Left_9323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_16_Left_9324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_16_Left_9325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_16_Left_9326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_16_Left_9327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_16_Left_9328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_16_Left_9329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_16_Left_9330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_16_Left_9331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_16_Left_9332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_16_Left_9333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_16_Left_9334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_16_Left_9335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_16_Left_9336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_16_Left_9337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_16_Left_9338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_16_Left_9339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_16_Left_9340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_16_Left_9341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_16_Left_9342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_16_Left_9343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_16_Left_9344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_16_Left_9345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_16_Left_9346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_16_Left_9347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_16_Left_9348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_16_Left_9349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_16_Left_9350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_16_Left_9351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_16_Left_9352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_16_Left_9353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_16_Left_9354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_16_Left_9355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_16_Left_9356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_16_Left_9357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_16_Left_9358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_16_Left_9359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_16_Left_9360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_16_Left_9361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_16_Left_9362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_16_Left_9363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_16_Left_9364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_16_Left_9365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_16_Left_9366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_16_Left_9367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_16_Left_9368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_16_Left_9369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_16_Left_9370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_16_Left_9371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_16_Left_9372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_16_Left_9373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_16_Left_9374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_16_Left_9375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_16_Left_9376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_16_Left_9377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_16_Left_9378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_16_Left_9379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_16_Left_9380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_16_Left_9381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_16_Left_9382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_16_Left_9383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_16_Left_9384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_16_Left_9385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_16_Left_9386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_16_Left_9387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_16_Left_9388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_16_Left_9389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_16_Left_9390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_16_Left_9391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_16_Left_9392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_16_Left_9393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_16_Left_9394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_16_Left_9395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_16_Right_9396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_16_Right_9397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_16_Right_9398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_16_Right_9399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_16_Right_9400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_16_Right_9401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_16_Right_9402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_16_Right_9403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_16_Right_9404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_16_Right_9405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_16_Right_9406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_16_Right_9407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_16_Right_9408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_16_Right_9409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_16_Right_9410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_16_Right_9411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_16_Right_9412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_16_Right_9413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_16_Right_9414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_16_Right_9415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_16_Right_9416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_16_Right_9417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_16_Right_9418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_16_Right_9419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_16_Right_9420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_16_Right_9421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_16_Right_9422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_16_Right_9423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_16_Right_9424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_16_Right_9425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_16_Right_9426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_16_Right_9427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_16_Right_9428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_16_Right_9429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_16_Right_9430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_16_Right_9431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_16_Right_9432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_16_Right_9433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_16_Right_9434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_16_Right_9435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_16_Right_9436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_16_Right_9437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_16_Right_9438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_16_Right_9439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_16_Right_9440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_16_Right_9441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_16_Right_9442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_16_Right_9443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_16_Right_9444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_16_Right_9445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_16_Right_9446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_16_Right_9447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_16_Right_9448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_16_Right_9449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_16_Right_9450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_16_Right_9451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_16_Right_9452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_16_Right_9453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_16_Right_9454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_16_Right_9455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_16_Right_9456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_16_Right_9457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_16_Right_9458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_16_Right_9459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_16_Right_9460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_16_Right_9461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_16_Right_9462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_16_Right_9463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_16_Right_9464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_16_Right_9465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_16_Right_9466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_16_Right_9467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_16_Right_9468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_16_Right_9469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_16_Right_9470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_16_Right_9471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_16_Right_9472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_16_Right_9473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_16_Right_9474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_16_Right_9475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_16_Right_9476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_16_Right_9477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_16_Right_9478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_16_Right_9479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_16_Right_9480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_16_Right_9481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_16_Right_9482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_16_Right_9483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_16_Right_9484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_16_Right_9485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_16_Right_9486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_16_Right_9487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_16_Right_9488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_16_Right_9489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_16_Right_9490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_16_Right_9491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_16_Right_9492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_16_Right_9493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_16_Right_9494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_16_Right_9495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_16_Right_9496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_16_Right_9497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_16_Right_9498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_16_Right_9499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_16_Right_9500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_16_Right_9501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_16_Right_9502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_16_Right_9503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_16_Right_9504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_16_Right_9505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_16_Right_9506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_16_Right_9507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_16_Right_9508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_16_Right_9509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_16_Right_9510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_16_Right_9511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_16_Right_9512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_16_Right_9513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_16_Right_9514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_16_Right_9515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_16_Right_9516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_16_Right_9517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_16_Right_9518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_16_Right_9519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_16_Right_9520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_16_Right_9521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_16_Right_9522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_16_Right_9523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_16_Right_9524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_16_Right_9525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_16_Right_9526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_16_Right_9527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_16_Right_9528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_16_Right_9529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_16_Right_9530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_16_Right_9531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_16_Right_9532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_16_Right_9533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_16_Right_9534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_16_Right_9535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_16_Right_9536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_16_Right_9537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_16_Right_9538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_16_Right_9539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_16_Right_9540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_16_Right_9541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_16_Right_9542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_16_Right_9543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_16_Right_9544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_16_Right_9545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_16_Right_9546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_16_Right_9547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_16_Right_9548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_16_Right_9549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_16_Right_9550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_16_Right_9551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_16_Right_9552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_16_Right_9553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_16_Right_9554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_16_Right_9555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_16_Right_9556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_16_Right_9557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_16_Right_9558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_16_Right_9559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_16_Right_9560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_16_Right_9561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_16_Right_9562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_16_Right_9563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_16_Right_9564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_16_Right_9565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_16_Right_9566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_16_Right_9567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_16_Right_9568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_16_Right_9569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_16_Right_9570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_16_Right_9571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_16_Right_9572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_16_Right_9573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_16_Right_9574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_16_Right_9575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_16_Right_9576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_16_Right_9577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_16_Right_9578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_16_Right_9579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_16_Right_9580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_16_Right_9581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_16_Right_9582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_16_Right_9583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_16_Right_9584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_16_Right_9585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_16_Right_9586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_16_Right_9587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_16_Right_9588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_16_Right_9589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_16_Right_9590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_16_Right_9591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_16_Right_9592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_16_Right_9593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_16_Right_9594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_16_Right_9595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_16_Right_9596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_16_Right_9597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_16_Right_9598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_16_Right_9599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_16_Right_9600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_16_Right_9601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_16_Right_9602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_16_Right_9603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_16_Right_9604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_16_Right_9605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_16_Right_9606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_16_Right_9607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_16_Right_9608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_16_Right_9609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_16_Right_9610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_16_Right_9611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_16_Right_9612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_16_Right_9613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_16_Right_9614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_16_Right_9615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_16_Right_9616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_16_Right_9617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_16_Right_9618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_16_Right_9619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_16_Right_9620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_16_Right_9621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_16_Right_9622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_16_Right_9623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_16_Right_9624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_16_Right_9625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_16_Right_9626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_16_Right_9627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_16_Right_9628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_16_Right_9629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_16_Right_9630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_16_Right_9631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_16_Right_9632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_16_Right_9633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_16_Right_9634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_16_Right_9635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_16_Right_9636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_16_Right_9637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_16_Right_9638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_16_Right_9639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_16_Right_9640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_16_Right_9641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_16_Right_9642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_16_Right_9643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_16_Right_9644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_16_Right_9645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_16_Right_9646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_16_Right_9647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_16_Right_9648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_16_Right_9649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_16_Right_9650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_16_Right_9651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_16_Right_9652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_16_Right_9653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_16_Right_9654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_16_Right_9655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_16_Right_9656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_16_Right_9657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_16_Right_9658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_16_Right_9659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_16_Right_9660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_16_Right_9661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_16_Right_9662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_16_Right_9663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_16_Right_9664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_16_Right_9665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_16_Right_9666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_16_Right_9667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_16_Right_9668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_16_Right_9669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_16_Right_9670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_16_Right_9671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_16_Right_9672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_16_Right_9673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_16_Right_9674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_16_Right_9675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_16_Right_9676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_16_Right_9677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_16_Right_9678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_16_Right_9679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_16_Right_9680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_16_Right_9681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_16_Right_9682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_16_Right_9683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_16_Right_9684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_16_Right_9685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_16_Right_9686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_16_Right_9687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_16_Right_9688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_16_Right_9689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_16_Right_9690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_16_Right_9691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_16_Right_9692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_16_Right_9693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_16_Right_9694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_16_Right_9695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_16_Right_9696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_16_Right_9697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_16_Right_9698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_16_Right_9699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_16_Right_9700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_16_Right_9701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_16_Right_9702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_16_Right_9703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_16_Right_9704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_16_Right_9705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_16_Right_9706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_16_Right_9707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_16_Right_9708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_16_Right_9709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_16_Right_9710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_16_Right_9711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_16_Right_9712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_16_Right_9713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_16_Right_9714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_16_Right_9715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_16_Right_9716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_16_Right_9717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_16_Right_9718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_16_Right_9719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_17_Left_9720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_17_Left_9721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_17_Left_9722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_17_Left_9723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_17_Left_9724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_17_Left_9725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_17_Left_9726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_17_Left_9727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_17_Left_9728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_17_Left_9729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_17_Left_9730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_17_Left_9731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_17_Left_9732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_17_Left_9733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_17_Left_9734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_17_Left_9735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_17_Left_9736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_17_Left_9737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_17_Left_9738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_17_Left_9739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_17_Left_9740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_17_Left_9741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_17_Left_9742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_17_Left_9743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_17_Left_9744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_17_Left_9745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_17_Left_9746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_17_Left_9747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_17_Left_9748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_17_Left_9749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_17_Left_9750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_17_Left_9751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_17_Left_9752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_17_Left_9753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_17_Left_9754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_17_Left_9755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_17_Left_9756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_17_Left_9757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_17_Left_9758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_17_Left_9759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_17_Left_9760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_17_Left_9761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_17_Left_9762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_17_Left_9763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_17_Left_9764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_17_Left_9765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_17_Left_9766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_17_Left_9767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_17_Left_9768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_17_Left_9769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_17_Left_9770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_17_Left_9771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_17_Left_9772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_17_Left_9773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_17_Left_9774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_17_Left_9775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_17_Left_9776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_17_Left_9777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_17_Left_9778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_17_Left_9779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_17_Left_9780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_17_Left_9781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_17_Left_9782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_17_Left_9783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_17_Left_9784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_17_Left_9785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_17_Left_9786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_17_Left_9787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_17_Left_9788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_17_Left_9789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_17_Left_9790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_17_Left_9791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_17_Left_9792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_17_Left_9793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_17_Left_9794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_17_Left_9795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_17_Left_9796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_17_Left_9797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_17_Left_9798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_17_Left_9799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_17_Left_9800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_17_Left_9801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_17_Left_9802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_17_Left_9803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_17_Left_9804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_17_Left_9805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_17_Left_9806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_17_Left_9807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_17_Left_9808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_17_Left_9809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_17_Left_9810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_17_Left_9811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_17_Left_9812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_17_Left_9813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_17_Left_9814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_17_Left_9815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_17_Left_9816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_17_Left_9817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_17_Left_9818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_17_Left_9819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_17_Left_9820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_17_Left_9821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_17_Left_9822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_17_Left_9823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_17_Left_9824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_17_Left_9825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_17_Left_9826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_17_Left_9827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_17_Left_9828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_17_Left_9829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_17_Left_9830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_17_Left_9831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_17_Left_9832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_17_Left_9833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_17_Left_9834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_17_Left_9835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_17_Left_9836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_17_Left_9837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_17_Left_9838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_17_Left_9839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_17_Left_9840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_17_Left_9841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_17_Left_9842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_17_Left_9843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_17_Left_9844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_17_Left_9845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_17_Left_9846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_17_Left_9847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_17_Left_9848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_17_Left_9849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_17_Left_9850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_17_Left_9851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_17_Left_9852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_17_Left_9853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_17_Left_9854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_17_Left_9855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_17_Left_9856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_17_Left_9857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_17_Left_9858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_17_Left_9859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_17_Left_9860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_17_Left_9861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_17_Left_9862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_17_Left_9863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_17_Left_9864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_17_Left_9865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_17_Left_9866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_17_Left_9867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_17_Left_9868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_17_Left_9869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_17_Left_9870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_17_Left_9871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_17_Left_9872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_17_Left_9873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_17_Left_9874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_17_Left_9875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_17_Left_9876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_17_Left_9877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_17_Left_9878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_17_Left_9879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_17_Left_9880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_17_Left_9881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_17_Left_9882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_17_Left_9883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_17_Left_9884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_17_Left_9885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_17_Left_9886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_17_Left_9887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_17_Left_9888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_17_Left_9889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_17_Left_9890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_17_Left_9891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_17_Left_9892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_17_Left_9893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_17_Left_9894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_17_Left_9895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_17_Left_9896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_17_Left_9897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_17_Left_9898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_17_Left_9899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_17_Left_9900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_17_Left_9901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_17_Left_9902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_17_Left_9903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_17_Left_9904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_17_Left_9905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_17_Left_9906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_17_Left_9907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_17_Left_9908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_17_Left_9909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_17_Left_9910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_17_Left_9911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_17_Left_9912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_17_Left_9913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_17_Left_9914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_17_Left_9915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_17_Left_9916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_17_Left_9917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_17_Left_9918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_17_Left_9919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_17_Left_9920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_17_Left_9921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_17_Left_9922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_17_Left_9923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_17_Left_9924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_17_Left_9925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_17_Left_9926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_17_Left_9927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_17_Left_9928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_17_Left_9929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_17_Left_9930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_17_Left_9931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_17_Left_9932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_17_Left_9933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_17_Left_9934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_17_Left_9935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_17_Left_9936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_17_Left_9937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_17_Left_9938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_17_Left_9939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_17_Left_9940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_17_Left_9941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_17_Left_9942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_17_Left_9943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_17_Left_9944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_17_Left_9945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_17_Left_9946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_17_Left_9947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_17_Left_9948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_17_Left_9949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_17_Left_9950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_17_Left_9951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_17_Left_9952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_17_Left_9953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_17_Left_9954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_17_Left_9955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_17_Left_9956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_17_Left_9957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_17_Left_9958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_17_Left_9959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_17_Left_9960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_17_Left_9961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_17_Left_9962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_17_Left_9963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_17_Left_9964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_17_Left_9965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_17_Left_9966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_17_Left_9967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_17_Left_9968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_17_Left_9969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_17_Left_9970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_17_Left_9971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_17_Left_9972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_17_Left_9973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_17_Left_9974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_17_Left_9975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_17_Left_9976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_17_Left_9977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_17_Left_9978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_17_Left_9979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_17_Left_9980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_17_Left_9981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_17_Left_9982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_17_Left_9983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_17_Left_9984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_17_Left_9985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_17_Left_9986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_17_Left_9987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_17_Left_9988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_17_Left_9989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_17_Left_9990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_17_Left_9991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_17_Left_9992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_17_Left_9993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_17_Left_9994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_17_Left_9995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_17_Left_9996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_17_Left_9997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_17_Left_9998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_17_Left_9999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_17_Left_10000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_17_Left_10001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_17_Left_10002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_17_Left_10003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_17_Left_10004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_17_Left_10005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_17_Left_10006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_17_Left_10007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_17_Left_10008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_17_Left_10009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_17_Left_10010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_17_Left_10011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_17_Left_10012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_17_Left_10013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_17_Left_10014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_17_Left_10015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_17_Left_10016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_17_Left_10017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_17_Left_10018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_17_Left_10019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_17_Left_10020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_17_Left_10021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_17_Left_10022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_17_Left_10023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_17_Left_10024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_17_Left_10025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_17_Left_10026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_17_Left_10027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_17_Left_10028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_17_Left_10029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_17_Left_10030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_17_Left_10031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_17_Left_10032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_17_Left_10033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_17_Left_10034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_17_Left_10035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_17_Left_10036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_17_Left_10037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_17_Left_10038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_17_Left_10039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_17_Left_10040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_17_Left_10041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_17_Left_10042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_17_Left_10043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Right_10044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Right_10045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Right_10046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Right_10047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_17_Right_10048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_17_Right_10049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_17_Right_10050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_17_Right_10051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_17_Right_10052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_17_Right_10053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_17_Right_10054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_17_Right_10055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_17_Right_10056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_17_Right_10057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_17_Right_10058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_17_Right_10059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_17_Right_10060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_17_Right_10061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_17_Right_10062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_17_Right_10063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_17_Right_10064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_17_Right_10065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_17_Right_10066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_17_Right_10067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_17_Right_10068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_17_Right_10069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_17_Right_10070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_17_Right_10071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_17_Right_10072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_17_Right_10073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_17_Right_10074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_17_Right_10075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_17_Right_10076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_17_Right_10077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_17_Right_10078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_17_Right_10079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_17_Right_10080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_17_Right_10081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_17_Right_10082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_17_Right_10083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_17_Right_10084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_17_Right_10085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_17_Right_10086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_17_Right_10087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_17_Right_10088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_17_Right_10089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_17_Right_10090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_17_Right_10091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_17_Right_10092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_17_Right_10093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_17_Right_10094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_17_Right_10095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_17_Right_10096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_17_Right_10097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_17_Right_10098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_17_Right_10099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_17_Right_10100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_17_Right_10101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_17_Right_10102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_17_Right_10103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_17_Right_10104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_17_Right_10105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_17_Right_10106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_17_Right_10107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_17_Right_10108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_17_Right_10109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_17_Right_10110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_17_Right_10111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_17_Right_10112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_17_Right_10113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_17_Right_10114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_17_Right_10115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_17_Right_10116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_17_Right_10117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_17_Right_10118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_17_Right_10119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_17_Right_10120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_17_Right_10121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_17_Right_10122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_17_Right_10123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_17_Right_10124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_17_Right_10125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_17_Right_10126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_17_Right_10127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_17_Right_10128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_17_Right_10129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_17_Right_10130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_17_Right_10131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_17_Right_10132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_17_Right_10133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_17_Right_10134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_17_Right_10135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_17_Right_10136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_17_Right_10137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_17_Right_10138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_17_Right_10139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_17_Right_10140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_17_Right_10141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_17_Right_10142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_17_Right_10143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_17_Right_10144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_17_Right_10145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_17_Right_10146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_17_Right_10147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_17_Right_10148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_17_Right_10149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_17_Right_10150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_17_Right_10151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_17_Right_10152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_17_Right_10153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_17_Right_10154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_17_Right_10155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_17_Right_10156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_17_Right_10157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_17_Right_10158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_17_Right_10159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_17_Right_10160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_17_Right_10161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_17_Right_10162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_17_Right_10163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_17_Right_10164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_17_Right_10165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_17_Right_10166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_17_Right_10167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_17_Right_10168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_17_Right_10169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_17_Right_10170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_17_Right_10171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_17_Right_10172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_17_Right_10173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_17_Right_10174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_17_Right_10175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_17_Right_10176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_17_Right_10177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_17_Right_10178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_17_Right_10179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_17_Right_10180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_17_Right_10181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_17_Right_10182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_17_Right_10183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_17_Right_10184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_17_Right_10185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_17_Right_10186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_17_Right_10187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_17_Right_10188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_17_Right_10189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_17_Right_10190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_17_Right_10191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_17_Right_10192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_17_Right_10193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_17_Right_10194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_17_Right_10195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_17_Right_10196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_17_Right_10197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_17_Right_10198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_17_Right_10199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_17_Right_10200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_17_Right_10201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_17_Right_10202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_17_Right_10203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_17_Right_10204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_17_Right_10205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_17_Right_10206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_17_Right_10207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_17_Right_10208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_17_Right_10209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_17_Right_10210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_17_Right_10211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_17_Right_10212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_17_Right_10213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_17_Right_10214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_17_Right_10215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_17_Right_10216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_17_Right_10217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_17_Right_10218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_17_Right_10219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_17_Right_10220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_17_Right_10221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_17_Right_10222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_17_Right_10223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_17_Right_10224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_17_Right_10225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_17_Right_10226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_17_Right_10227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_17_Right_10228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_17_Right_10229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_17_Right_10230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_17_Right_10231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_17_Right_10232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_17_Right_10233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_17_Right_10234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_17_Right_10235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_17_Right_10236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_17_Right_10237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_17_Right_10238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_17_Right_10239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_17_Right_10240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_17_Right_10241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_17_Right_10242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_17_Right_10243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_17_Right_10244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_17_Right_10245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_17_Right_10246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_17_Right_10247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_17_Right_10248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_17_Right_10249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_17_Right_10250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_17_Right_10251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_17_Right_10252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_17_Right_10253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_17_Right_10254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_17_Right_10255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_17_Right_10256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_17_Right_10257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_17_Right_10258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_17_Right_10259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_17_Right_10260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_17_Right_10261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_17_Right_10262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_17_Right_10263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_17_Right_10264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_17_Right_10265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_17_Right_10266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_17_Right_10267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_17_Right_10268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_17_Right_10269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_17_Right_10270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_17_Right_10271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_17_Right_10272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_17_Right_10273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_17_Right_10274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_17_Right_10275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_17_Right_10276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_17_Right_10277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_17_Right_10278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_17_Right_10279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_17_Right_10280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_17_Right_10281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_17_Right_10282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_17_Right_10283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_17_Right_10284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_17_Right_10285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_17_Right_10286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_17_Right_10287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_17_Right_10288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_17_Right_10289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_17_Right_10290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_17_Right_10291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_17_Right_10292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_17_Right_10293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_17_Right_10294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_17_Right_10295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_17_Right_10296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_17_Right_10297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_17_Right_10298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_17_Right_10299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_17_Right_10300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_17_Right_10301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_17_Right_10302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_17_Right_10303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_17_Right_10304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_17_Right_10305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_17_Right_10306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_17_Right_10307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_17_Right_10308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_17_Right_10309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_17_Right_10310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_17_Right_10311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_17_Right_10312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_17_Right_10313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_17_Right_10314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_17_Right_10315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_17_Right_10316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_17_Right_10317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_17_Right_10318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_17_Right_10319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_17_Right_10320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_17_Right_10321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_17_Right_10322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_17_Right_10323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_17_Right_10324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_17_Right_10325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_17_Right_10326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_17_Right_10327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_17_Right_10328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_17_Right_10329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_17_Right_10330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_17_Right_10331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_17_Right_10332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_17_Right_10333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_17_Right_10334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_17_Right_10335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_17_Right_10336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_17_Right_10337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_17_Right_10338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_17_Right_10339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_17_Right_10340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_17_Right_10341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_17_Right_10342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_17_Right_10343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_17_Right_10344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_17_Right_10345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_17_Right_10346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_17_Right_10347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_17_Right_10348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_17_Right_10349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_17_Right_10350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_17_Right_10351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_17_Right_10352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_17_Right_10353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_17_Right_10354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_17_Right_10355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_17_Right_10356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_17_Right_10357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_17_Right_10358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_17_Right_10359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_17_Right_10360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_17_Right_10361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_17_Right_10362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_17_Right_10363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_17_Right_10364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_17_Right_10365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_17_Right_10366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_17_Right_10367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_17_Right_10368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_17_Right_10369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_17_Right_10370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_17_Right_10371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Left_10372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Left_10373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Left_10374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Left_10375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_2_10376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_2_10377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_2_10378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_2_10379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_2_10380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_2_10381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_2_10382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_2_10383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_10384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_10385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_10386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_10387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_10388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_10389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_10390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_10391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_10392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_10393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_10394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_10395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_10396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_10397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_10398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_10399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_10400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_10401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_10402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_10403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_10404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_10405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_10406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_10407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_10408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_10409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_10410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_10411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_10412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_10413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_10414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_10415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_10416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2_10417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2_10418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2_10419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2_10420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2_10421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2_10422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2_10423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2_10424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2_10425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2_10426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2_10427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2_10428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2_10429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2_10430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2_10431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2_10432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2_10433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2_10434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2_10435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2_10436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2_10437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2_10438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2_10439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2_10440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2_10441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2_10442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2_10443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2_10444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2_10445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2_10446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2_10447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2_10448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2_10449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2_10450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2_10451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2_10452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2_10453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2_10454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2_10455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2_10456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2_10457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2_10458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2_10459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2_10460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2_10461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2_10462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2_10463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2_10464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2_10465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2_10466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2_10467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2_10468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2_10469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2_10470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2_10471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2_10472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2_10473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2_10474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2_10475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2_10476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2_10477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2_10478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2_10479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2_10480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2_10481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2_10482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2_10483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_2_10484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_2_10485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_2_10486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_2_10487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_2_10488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_2_10489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_2_10490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_2_10491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_2_10492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_2_10493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_2_10494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_2_10495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_2_10496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_2_10497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_2_10498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_2_10499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_2_10500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_2_10501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_2_10502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_2_10503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_2_10504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_2_10505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_2_10506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_2_10507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_2_10508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_2_10509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_2_10510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_2_10511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_2_10512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_2_10513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_2_10514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_2_10515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_2_10516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_2_10517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_2_10518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_2_10519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_2_10520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_2_10521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_2_10522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_2_10523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_2_10524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_2_10525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_2_10526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_2_10527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_2_10528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_2_10529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_2_10530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_2_10531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_2_10532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_2_10533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_2_10534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_2_10535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_2_10536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_10684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_10756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_10828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_10976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_2_10977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_3_10978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_4_10979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_5_10980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_6_10981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_7_10982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_8_10983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_9_10984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_10_10985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_11_10986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_12_10987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_13_10988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_14_10989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_15_10990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_16_10991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_3_10992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_4_10993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_5_10994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_6_10995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_7_10996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_8_10997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_9_10998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_10_10999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_11_11000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_12_11001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_13_11002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_14_11003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_15_11004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_16_11005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_3_11006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_4_11007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_5_11008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_6_11009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_7_11010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_8_11011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_9_11012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_10_11013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_11_11014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_12_11015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_13_11016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_14_11017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_15_11018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_16_11019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_3_11020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_4_11021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_5_11022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_6_11023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_7_11024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_8_11025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_9_11026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_10_11027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_11_11028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_12_11029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_13_11030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_14_11031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_15_11032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_16_11033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_3_11034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_4_11035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_5_11036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_6_11037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_7_11038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_8_11039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_9_11040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_10_11041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_11_11042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_12_11043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_13_11044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_14_11045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_15_11046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_16_11047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_3_11048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_4_11049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_5_11050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_6_11051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_7_11052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_8_11053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_9_11054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_10_11055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_11_11056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_12_11057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_13_11058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_14_11059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_15_11060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_16_11061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_3_11062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_4_11063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_5_11064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_6_11065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_7_11066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_8_11067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_9_11068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_10_11069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_11_11070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_12_11071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_13_11072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_14_11073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_15_11074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_16_11075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_3_11076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_4_11077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_5_11078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_6_11079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_7_11080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_8_11081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_9_11082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_10_11083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_11_11084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_12_11085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_13_11086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_14_11087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_15_11088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_16_11089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_3_11090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_4_11091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_5_11092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_6_11093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_7_11094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_8_11095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_9_11096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_10_11097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_11_11098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_12_11099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_13_11100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_14_11101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_15_11102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_16_11103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_3_11104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_4_11105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_5_11106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_6_11107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_7_11108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_8_11109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_9_11110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_10_11111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_11_11112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_12_11113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_13_11114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_14_11115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_15_11116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_16_11117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_3_11118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_4_11119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_5_11120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_6_11121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_7_11122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_8_11123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_9_11124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_10_11125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_11_11126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_12_11127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_13_11128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_14_11129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_15_11130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_16_11131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_3_11132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_4_11133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_5_11134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_6_11135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_7_11136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_8_11137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_9_11138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_10_11139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_11_11140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_12_11141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_13_11142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_14_11143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_15_11144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_16_11145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_3_11146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_4_11147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_5_11148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_6_11149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_7_11150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_8_11151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_9_11152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_10_11153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_11_11154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_12_11155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_13_11156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_14_11157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_15_11158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_16_11159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_3_11160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_4_11161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_5_11162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_6_11163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_7_11164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_8_11165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_9_11166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_10_11167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_11_11168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_12_11169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_13_11170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_14_11171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_15_11172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_16_11173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_3_11174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_4_11175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_5_11176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_6_11177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_7_11178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_8_11179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_9_11180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_10_11181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_11_11182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_12_11183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_13_11184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_14_11185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_15_11186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_16_11187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_3_11188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_4_11189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_5_11190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_6_11191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_7_11192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_8_11193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_9_11194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_10_11195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_11_11196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_12_11197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_13_11198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_14_11199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_15_11200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_16_11201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_3_11202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_4_11203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_5_11204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_6_11205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_7_11206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_8_11207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_9_11208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_10_11209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_11_11210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_12_11211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_13_11212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_14_11213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_15_11214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_16_11215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_3_11216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_4_11217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_5_11218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_6_11219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_7_11220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_8_11221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_9_11222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_10_11223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_11_11224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_12_11225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_13_11226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_14_11227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_15_11228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_16_11229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_3_11230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_4_11231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_5_11232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_6_11233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_7_11234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_8_11235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_9_11236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_10_11237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_11_11238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_12_11239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_13_11240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_14_11241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_15_11242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_16_11243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_3_11244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_4_11245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_5_11246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_6_11247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_7_11248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_8_11249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_9_11250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_10_11251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_11_11252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_12_11253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_13_11254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_14_11255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_15_11256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_16_11257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_3_11258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_4_11259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_5_11260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_6_11261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_7_11262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_8_11263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_9_11264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_10_11265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_11_11266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_12_11267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_13_11268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_14_11269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_15_11270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_16_11271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_3_11272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_4_11273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_5_11274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_6_11275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_7_11276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_8_11277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_9_11278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_10_11279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_11_11280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_12_11281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_13_11282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_14_11283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_15_11284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_16_11285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_3_11286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_4_11287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_5_11288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_6_11289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_7_11290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_8_11291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_9_11292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_10_11293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_11_11294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_12_11295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_13_11296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_14_11297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_15_11298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_16_11299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_3_11300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_4_11301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_5_11302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_6_11303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_7_11304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_8_11305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_9_11306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_10_11307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_11_11308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_12_11309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_13_11310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_14_11311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_15_11312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_16_11313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_3_11314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_4_11315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_5_11316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_6_11317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_7_11318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_8_11319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_9_11320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_10_11321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_11_11322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_12_11323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_13_11324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_14_11325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_15_11326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_16_11327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_3_11328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_4_11329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_5_11330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_6_11331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_7_11332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_8_11333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_9_11334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_10_11335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_11_11336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_12_11337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_13_11338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_14_11339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_15_11340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_16_11341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_3_11342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_4_11343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_5_11344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_6_11345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_7_11346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_8_11347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_9_11348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_10_11349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_11_11350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_12_11351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_13_11352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_14_11353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_15_11354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_16_11355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_3_11356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_4_11357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_5_11358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_6_11359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_7_11360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_8_11361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_9_11362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_10_11363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_11_11364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_12_11365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_13_11366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_14_11367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_15_11368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_16_11369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_3_11370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_4_11371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_5_11372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_6_11373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_7_11374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_8_11375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_9_11376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_10_11377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_11_11378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_12_11379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_13_11380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_14_11381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_15_11382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_16_11383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_3_11384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_4_11385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_5_11386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_6_11387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_7_11388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_8_11389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_9_11390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_10_11391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_11_11392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_12_11393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_13_11394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_14_11395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_15_11396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_16_11397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_3_11398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_4_11399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_5_11400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_6_11401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_7_11402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_8_11403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_9_11404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_10_11405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_11_11406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_12_11407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_13_11408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_14_11409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_15_11410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_16_11411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_3_11412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_4_11413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_5_11414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_6_11415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_7_11416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_8_11417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_9_11418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_10_11419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_11_11420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_12_11421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_13_11422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_14_11423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_15_11424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_16_11425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_3_11426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_4_11427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_5_11428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_6_11429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_7_11430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_8_11431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_9_11432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_10_11433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_11_11434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_12_11435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_13_11436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_14_11437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_15_11438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_16_11439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_3_11440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_4_11441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_5_11442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_6_11443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_7_11444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_8_11445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_9_11446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_10_11447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_11_11448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_12_11449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_13_11450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_14_11451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_15_11452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_16_11453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_3_11454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_4_11455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_5_11456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_6_11457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_7_11458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_8_11459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_9_11460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_10_11461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_11_11462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_12_11463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_13_11464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_14_11465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_15_11466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_16_11467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_3_11468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_4_11469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_5_11470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_6_11471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_7_11472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_8_11473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_9_11474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_10_11475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_11_11476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_12_11477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_13_11478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_14_11479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_15_11480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_16_11481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_3_11482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_4_11483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_5_11484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_6_11485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_7_11486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_8_11487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_9_11488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_10_11489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_11_11490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_12_11491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_13_11492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_14_11493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_15_11494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_16_11495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_3_11496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_4_11497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_5_11498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_6_11499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_7_11500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_8_11501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_9_11502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_10_11503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_11_11504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_12_11505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_13_11506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_14_11507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_15_11508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_16_11509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_3_11510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_4_11511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_5_11512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_6_11513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_7_11514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_8_11515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_9_11516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_10_11517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_11_11518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_12_11519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_13_11520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_14_11521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_15_11522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_16_11523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_3_11524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_4_11525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_5_11526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_6_11527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_7_11528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_8_11529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_9_11530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_10_11531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_11_11532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_12_11533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_13_11534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_14_11535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_15_11536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_16_11537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_3_11538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_4_11539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_5_11540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_6_11541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_7_11542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_8_11543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_9_11544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_10_11545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_11_11546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_12_11547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_13_11548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_14_11549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_15_11550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_16_11551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_3_11552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_4_11553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_5_11554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_6_11555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_7_11556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_8_11557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_9_11558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_10_11559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_11_11560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_12_11561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_13_11562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_14_11563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_15_11564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_16_11565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_3_11566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_4_11567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_5_11568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_6_11569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_7_11570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_8_11571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_9_11572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_10_11573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_11_11574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_12_11575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_13_11576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_14_11577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_15_11578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_16_11579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_3_11580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_4_11581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_5_11582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_6_11583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_7_11584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_8_11585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_9_11586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_10_11587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_11_11588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_12_11589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_13_11590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_14_11591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_15_11592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_16_11593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_3_11594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_4_11595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_5_11596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_6_11597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_7_11598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_8_11599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_9_11600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_10_11601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_11_11602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_12_11603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_13_11604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_14_11605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_15_11606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_16_11607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_3_11608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_4_11609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_5_11610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_6_11611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_7_11612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_8_11613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_9_11614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_10_11615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_11_11616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_12_11617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_13_11618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_14_11619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_15_11620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_16_11621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_3_11622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_4_11623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_5_11624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_6_11625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_7_11626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_8_11627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_9_11628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_10_11629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_11_11630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_12_11631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_13_11632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_14_11633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_15_11634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_16_11635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3_11636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_4_11637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_5_11638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_6_11639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_7_11640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_8_11641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_9_11642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_10_11643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_11_11644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_12_11645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_13_11646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_14_11647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_15_11648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_16_11649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3_11650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_4_11651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_5_11652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_6_11653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_7_11654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_8_11655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_9_11656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_10_11657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_11_11658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_12_11659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_13_11660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_14_11661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_15_11662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_16_11663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3_11664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_4_11665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_5_11666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_6_11667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_7_11668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_8_11669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_9_11670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_10_11671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_11_11672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_12_11673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_13_11674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_14_11675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_15_11676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_16_11677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3_11678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_4_11679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_5_11680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_6_11681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_7_11682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_8_11683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_9_11684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_10_11685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_11_11686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_12_11687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_13_11688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_14_11689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_15_11690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_16_11691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3_11692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_4_11693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_5_11694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_6_11695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_7_11696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_8_11697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_9_11698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_10_11699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_11_11700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_12_11701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_13_11702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_14_11703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_15_11704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_16_11705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3_11706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_4_11707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_5_11708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_6_11709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_7_11710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_8_11711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_9_11712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_10_11713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_11_11714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_12_11715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_13_11716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_14_11717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_15_11718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_16_11719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3_11720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_4_11721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_5_11722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_6_11723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_7_11724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_8_11725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_9_11726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_10_11727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_11_11728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_12_11729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_13_11730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_14_11731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_15_11732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_16_11733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3_11734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_4_11735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_5_11736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_6_11737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_7_11738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_8_11739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_9_11740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_10_11741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_11_11742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_12_11743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_13_11744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_14_11745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_15_11746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_16_11747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3_11748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_4_11749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_5_11750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_6_11751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_7_11752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_8_11753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_9_11754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_10_11755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_11_11756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_12_11757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_13_11758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_14_11759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_15_11760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_16_11761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3_11762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_4_11763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_5_11764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_6_11765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_7_11766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_8_11767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_9_11768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_10_11769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_11_11770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_12_11771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_13_11772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_14_11773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_15_11774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_16_11775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3_11776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_4_11777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_5_11778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_6_11779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_7_11780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_8_11781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_9_11782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_10_11783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_11_11784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_12_11785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_13_11786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_14_11787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_15_11788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_16_11789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3_11790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_4_11791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_5_11792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_6_11793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_7_11794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_8_11795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_9_11796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_10_11797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_11_11798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_12_11799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_13_11800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_14_11801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_15_11802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_16_11803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3_11804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_4_11805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_5_11806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_6_11807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_7_11808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_8_11809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_9_11810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_10_11811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_11_11812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_12_11813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_13_11814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_14_11815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_15_11816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_16_11817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3_11818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_4_11819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_5_11820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_6_11821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_7_11822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_8_11823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_9_11824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_10_11825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_11_11826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_12_11827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_13_11828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_14_11829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_15_11830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_16_11831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3_11832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_4_11833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_5_11834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_6_11835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_7_11836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_8_11837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_9_11838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_10_11839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_11_11840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_12_11841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_13_11842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_14_11843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_15_11844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_16_11845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3_11846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_4_11847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_5_11848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_6_11849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_7_11850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_8_11851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_9_11852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_10_11853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_11_11854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_12_11855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_13_11856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_14_11857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_15_11858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_16_11859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3_11860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_4_11861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_5_11862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_6_11863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_7_11864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_8_11865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_9_11866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_10_11867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_11_11868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_12_11869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_13_11870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_14_11871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_15_11872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_16_11873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3_11874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_4_11875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_5_11876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_6_11877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_7_11878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_8_11879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_9_11880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_10_11881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_11_11882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_12_11883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_13_11884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_14_11885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_15_11886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_16_11887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3_11888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4_11889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_5_11890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_6_11891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_7_11892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_8_11893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_9_11894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_10_11895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_11_11896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_12_11897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_13_11898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_14_11899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_15_11900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_16_11901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3_11902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4_11903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_5_11904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_6_11905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_7_11906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_8_11907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_9_11908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_10_11909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_11_11910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_12_11911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_13_11912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_14_11913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_15_11914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_16_11915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3_11916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4_11917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_5_11918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_6_11919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_7_11920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_8_11921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_9_11922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_10_11923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_11_11924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_12_11925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_13_11926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_14_11927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_15_11928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_16_11929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3_11930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4_11931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_5_11932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_6_11933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_7_11934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_8_11935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_9_11936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_10_11937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_11_11938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_12_11939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_13_11940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_14_11941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_15_11942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_16_11943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3_11944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4_11945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_5_11946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_6_11947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_7_11948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_8_11949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_9_11950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_10_11951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_11_11952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_12_11953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_13_11954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_14_11955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_15_11956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_16_11957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3_11958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4_11959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_5_11960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_6_11961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_7_11962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_8_11963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_9_11964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_10_11965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_11_11966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_12_11967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_13_11968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_14_11969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_15_11970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_16_11971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3_11972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4_11973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_5_11974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_6_11975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_7_11976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_8_11977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_9_11978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_10_11979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_11_11980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_12_11981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_13_11982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_14_11983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_15_11984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_16_11985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3_11986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4_11987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_5_11988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_6_11989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_7_11990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_8_11991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_9_11992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_10_11993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_11_11994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_12_11995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_13_11996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_14_11997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_15_11998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_16_11999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3_12000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4_12001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_5_12002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_6_12003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_7_12004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_8_12005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_9_12006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_10_12007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_11_12008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_12_12009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_13_12010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_14_12011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_15_12012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_16_12013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3_12014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4_12015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_5_12016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_6_12017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_7_12018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_8_12019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_9_12020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_10_12021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_11_12022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_12_12023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_13_12024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_14_12025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_15_12026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_16_12027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3_12028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4_12029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_5_12030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_6_12031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_7_12032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_8_12033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_9_12034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_10_12035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_11_12036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_12_12037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_13_12038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_14_12039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_15_12040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_16_12041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3_12042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4_12043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_5_12044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_6_12045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_7_12046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_8_12047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_9_12048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_10_12049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_11_12050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_12_12051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_13_12052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_14_12053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_15_12054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_16_12055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3_12056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4_12057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_5_12058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_6_12059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_7_12060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_8_12061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_9_12062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_10_12063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_11_12064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_12_12065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_13_12066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_14_12067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_15_12068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_16_12069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3_12070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4_12071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_5_12072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_6_12073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_7_12074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_8_12075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_9_12076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_10_12077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_11_12078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_12_12079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_13_12080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_14_12081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_15_12082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_16_12083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3_12084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4_12085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_5_12086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_6_12087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_7_12088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_8_12089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_9_12090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_10_12091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_11_12092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_12_12093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_13_12094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_14_12095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_15_12096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_16_12097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3_12098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4_12099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_5_12100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_6_12101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_7_12102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_8_12103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_9_12104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_10_12105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_11_12106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_12_12107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_13_12108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_14_12109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_15_12110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_16_12111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3_12112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4_12113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_5_12114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_6_12115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_7_12116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_8_12117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_9_12118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_10_12119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_11_12120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_12_12121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_13_12122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_14_12123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_15_12124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_16_12125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3_12126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4_12127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_5_12128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_6_12129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_7_12130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_8_12131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_9_12132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_10_12133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_11_12134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_12_12135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_13_12136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_14_12137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_15_12138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_16_12139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3_12140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4_12141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5_12142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_6_12143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_7_12144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_8_12145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_9_12146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_10_12147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_11_12148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_12_12149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_13_12150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_14_12151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_15_12152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_16_12153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3_12154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4_12155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5_12156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_6_12157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_7_12158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_8_12159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_9_12160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_10_12161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_11_12162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_12_12163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_13_12164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_14_12165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_15_12166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_16_12167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3_12168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_4_12169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5_12170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_6_12171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_7_12172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_8_12173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_9_12174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_10_12175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_11_12176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_12_12177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_13_12178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_14_12179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_15_12180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_16_12181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3_12182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_4_12183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5_12184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_6_12185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_7_12186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_8_12187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_9_12188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_10_12189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_11_12190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_12_12191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_13_12192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_14_12193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_15_12194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_16_12195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3_12196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_4_12197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5_12198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_6_12199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_7_12200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_8_12201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_9_12202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_10_12203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_11_12204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_12_12205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_13_12206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_14_12207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_15_12208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_16_12209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3_12210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_4_12211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5_12212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_6_12213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_7_12214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_8_12215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_9_12216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_10_12217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_11_12218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_12_12219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_13_12220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_14_12221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_15_12222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_16_12223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3_12224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_4_12225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5_12226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_6_12227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_7_12228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_8_12229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_9_12230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_10_12231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_11_12232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_12_12233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_13_12234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_14_12235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_15_12236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_16_12237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3_12238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_4_12239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5_12240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_6_12241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_7_12242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_8_12243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_9_12244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_10_12245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_11_12246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_12_12247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_13_12248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_14_12249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_15_12250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_16_12251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3_12252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_4_12253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5_12254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_6_12255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_7_12256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_8_12257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_9_12258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_10_12259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_11_12260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_12_12261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_13_12262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_14_12263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_15_12264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_16_12265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_3_12266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_4_12267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5_12268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_6_12269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_7_12270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_8_12271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_9_12272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_10_12273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_11_12274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_12_12275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_13_12276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_14_12277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_15_12278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_16_12279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_3_12280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_4_12281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5_12282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_6_12283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_7_12284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_8_12285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_9_12286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_10_12287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_11_12288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_12_12289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_13_12290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_14_12291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_15_12292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_16_12293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_3_12294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_4_12295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5_12296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_6_12297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_7_12298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_8_12299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_9_12300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_10_12301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_11_12302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_12_12303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_13_12304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_14_12305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_15_12306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_16_12307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_3_12308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_4_12309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5_12310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_6_12311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_7_12312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_8_12313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_9_12314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_10_12315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_11_12316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_12_12317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_13_12318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_14_12319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_15_12320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_16_12321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_3_12322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_4_12323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5_12324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_6_12325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_7_12326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_8_12327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_9_12328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_10_12329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_11_12330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_12_12331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_13_12332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_14_12333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_15_12334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_16_12335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_3_12336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_4_12337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5_12338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_6_12339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_7_12340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_8_12341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_9_12342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_10_12343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_11_12344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_12_12345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_13_12346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_14_12347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_15_12348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_16_12349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_3_12350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_4_12351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_5_12352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_6_12353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_7_12354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_8_12355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_9_12356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_10_12357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_11_12358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_12_12359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_13_12360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_14_12361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_15_12362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_16_12363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_3_12364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_4_12365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_5_12366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_6_12367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_7_12368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_8_12369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_9_12370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_10_12371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_11_12372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_12_12373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_13_12374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_14_12375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_15_12376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_16_12377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_3_12378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_4_12379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_5_12380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_6_12381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_7_12382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_8_12383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_9_12384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_10_12385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_11_12386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_12_12387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_13_12388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_14_12389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_15_12390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_16_12391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_3_12392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_4_12393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_5_12394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_6_12395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_7_12396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_8_12397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_9_12398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_10_12399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_11_12400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_12_12401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_13_12402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_14_12403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_15_12404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_16_12405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_3_12406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_4_12407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_5_12408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_6_12409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_7_12410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_8_12411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_9_12412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_10_12413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_11_12414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_12_12415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_13_12416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_14_12417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_15_12418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_16_12419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_3_12420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_4_12421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_5_12422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_6_12423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_7_12424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_8_12425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_9_12426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_10_12427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_11_12428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_12_12429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_13_12430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_14_12431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_15_12432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_16_12433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_3_12434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_4_12435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_5_12436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_6_12437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_7_12438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_8_12439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_9_12440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_10_12441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_11_12442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_12_12443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_13_12444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_14_12445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_15_12446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_16_12447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_3_12448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_4_12449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_5_12450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_6_12451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_7_12452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_8_12453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_9_12454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_10_12455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_11_12456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_12_12457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_13_12458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_14_12459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_15_12460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_16_12461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_3_12462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_4_12463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_5_12464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_6_12465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_7_12466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_8_12467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_9_12468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_10_12469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_11_12470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_12_12471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_13_12472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_14_12473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_15_12474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_16_12475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_3_12476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_4_12477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_5_12478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_6_12479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_7_12480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_8_12481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_9_12482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_10_12483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_11_12484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_12_12485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_13_12486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_14_12487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_15_12488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_16_12489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_3_12490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_4_12491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_5_12492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_6_12493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_7_12494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_8_12495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_9_12496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_10_12497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_11_12498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_12_12499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_13_12500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_14_12501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_15_12502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_16_12503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3_12504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_4_12505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_5_12506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_6_12507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_7_12508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_8_12509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_9_12510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_10_12511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_11_12512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_12_12513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_13_12514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_14_12515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_15_12516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_16_12517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3_12518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_4_12519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_5_12520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_6_12521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_7_12522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_8_12523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_9_12524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_10_12525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_11_12526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_12_12527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_13_12528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_14_12529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_15_12530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_16_12531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3_12532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_4_12533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_5_12534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_6_12535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_7_12536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_8_12537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_9_12538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_10_12539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_11_12540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_12_12541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_13_12542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_14_12543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_15_12544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_16_12545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3_12546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_4_12547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_5_12548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_6_12549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_7_12550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_8_12551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_9_12552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_10_12553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_11_12554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_12_12555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_13_12556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_14_12557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_15_12558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_16_12559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3_12560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_4_12561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_5_12562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_6_12563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_7_12564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_8_12565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_9_12566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_10_12567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_11_12568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_12_12569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_13_12570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_14_12571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_15_12572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_16_12573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3_12574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_4_12575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_5_12576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_6_12577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_7_12578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_8_12579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_9_12580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_10_12581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_11_12582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_12_12583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_13_12584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_14_12585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_15_12586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_16_12587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3_12588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_4_12589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_5_12590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_6_12591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_7_12592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_8_12593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_9_12594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_10_12595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_11_12596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_12_12597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_13_12598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_14_12599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_15_12600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_16_12601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3_12602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_4_12603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_5_12604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_6_12605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_7_12606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_8_12607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_9_12608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_10_12609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_11_12610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_12_12611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_13_12612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_14_12613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_15_12614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_16_12615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3_12616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_4_12617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_5_12618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_6_12619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_7_12620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_8_12621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_9_12622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_10_12623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_11_12624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_12_12625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_13_12626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_14_12627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_15_12628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_16_12629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3_12630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_4_12631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_5_12632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_6_12633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_7_12634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_8_12635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_9_12636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_10_12637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_11_12638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_12_12639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_13_12640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_14_12641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_15_12642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_16_12643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3_12644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_4_12645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_5_12646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_6_12647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_7_12648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_8_12649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_9_12650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_10_12651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_11_12652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_12_12653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_13_12654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_14_12655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_15_12656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_16_12657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3_12658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_4_12659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_5_12660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_6_12661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_7_12662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_8_12663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_9_12664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_10_12665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_11_12666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_12_12667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_13_12668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_14_12669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_15_12670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_16_12671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3_12672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_4_12673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_5_12674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_6_12675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_7_12676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_8_12677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_9_12678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_10_12679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_11_12680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_12_12681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_13_12682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_14_12683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_15_12684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_16_12685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3_12686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_4_12687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_5_12688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_6_12689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_7_12690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_8_12691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_9_12692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_10_12693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_11_12694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_12_12695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_13_12696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_14_12697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_15_12698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_16_12699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3_12700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_4_12701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_5_12702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_6_12703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_7_12704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_8_12705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_9_12706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_10_12707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_11_12708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_12_12709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_13_12710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_14_12711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_15_12712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_16_12713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3_12714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_4_12715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_5_12716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_6_12717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_7_12718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_8_12719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_9_12720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_10_12721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_11_12722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_12_12723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_13_12724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_14_12725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_15_12726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_16_12727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3_12728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_4_12729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_5_12730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_6_12731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_7_12732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_8_12733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_9_12734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_10_12735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_11_12736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_12_12737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_13_12738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_14_12739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_15_12740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_16_12741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3_12742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_4_12743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_5_12744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_6_12745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_7_12746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_8_12747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_9_12748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_10_12749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_11_12750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_12_12751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_13_12752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_14_12753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_15_12754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_16_12755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3_12756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_4_12757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_5_12758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_6_12759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_7_12760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_8_12761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_9_12762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_10_12763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_11_12764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_12_12765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_13_12766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_14_12767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_15_12768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_16_12769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3_12770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_4_12771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_5_12772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_6_12773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_7_12774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_8_12775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_9_12776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_10_12777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_11_12778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_12_12779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_13_12780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_14_12781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_15_12782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_16_12783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3_12784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_4_12785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_5_12786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_6_12787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_7_12788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_8_12789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_9_12790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_10_12791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_11_12792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_12_12793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_13_12794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_14_12795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_15_12796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_16_12797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3_12798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_4_12799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_5_12800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_6_12801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_7_12802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_8_12803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_9_12804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_10_12805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_11_12806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_12_12807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_13_12808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_14_12809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_15_12810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_16_12811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3_12812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_4_12813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_5_12814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_6_12815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_7_12816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_8_12817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_9_12818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_10_12819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_11_12820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_12_12821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_13_12822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_14_12823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_15_12824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_16_12825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3_12826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_4_12827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_5_12828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_6_12829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_7_12830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_8_12831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_9_12832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_10_12833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_11_12834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_12_12835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_13_12836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_14_12837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_15_12838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_16_12839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3_12840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_4_12841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_5_12842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_6_12843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_7_12844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_8_12845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_9_12846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_10_12847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_11_12848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_12_12849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_13_12850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_14_12851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_15_12852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_16_12853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3_12854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_4_12855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_5_12856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_6_12857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_7_12858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_8_12859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_9_12860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_10_12861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_11_12862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_12_12863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_13_12864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_14_12865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_15_12866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_16_12867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3_12868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_4_12869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_5_12870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_6_12871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_7_12872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_8_12873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_9_12874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_10_12875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_11_12876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_12_12877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_13_12878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_14_12879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_15_12880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_16_12881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3_12882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_4_12883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_5_12884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_6_12885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_7_12886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_8_12887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_9_12888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_10_12889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_11_12890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_12_12891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_13_12892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_14_12893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_15_12894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_16_12895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3_12896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_4_12897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_5_12898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_6_12899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_7_12900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_8_12901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_9_12902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_10_12903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_11_12904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_12_12905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_13_12906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_14_12907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_15_12908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_16_12909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3_12910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_4_12911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_5_12912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_6_12913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_7_12914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_8_12915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_9_12916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_10_12917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_11_12918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_12_12919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_13_12920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_14_12921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_15_12922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_16_12923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3_12924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_4_12925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_5_12926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_6_12927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_7_12928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_8_12929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_9_12930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_10_12931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_11_12932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_12_12933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_13_12934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_14_12935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_15_12936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_16_12937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3_12938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_4_12939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_5_12940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_6_12941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_7_12942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_8_12943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_9_12944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_10_12945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_11_12946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_12_12947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_13_12948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_14_12949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_15_12950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_16_12951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3_12952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_4_12953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_5_12954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_6_12955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_7_12956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_8_12957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_9_12958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_10_12959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_11_12960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_12_12961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_13_12962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_14_12963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_15_12964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_16_12965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3_12966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_4_12967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_5_12968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_6_12969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_7_12970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_8_12971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_9_12972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_10_12973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_11_12974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_12_12975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_13_12976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_14_12977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_15_12978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_16_12979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3_12980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_4_12981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_5_12982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_6_12983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_7_12984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_8_12985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_9_12986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_10_12987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_11_12988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_12_12989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_13_12990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_14_12991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_15_12992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_16_12993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3_12994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_4_12995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_5_12996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_6_12997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_7_12998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_8_12999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_9_13000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_10_13001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_11_13002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_12_13003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_13_13004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_14_13005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_15_13006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_16_13007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3_13008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_4_13009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_5_13010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_6_13011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_7_13012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_8_13013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_9_13014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_10_13015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_11_13016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_12_13017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_13_13018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_14_13019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_15_13020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_16_13021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3_13022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_4_13023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_5_13024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_6_13025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_7_13026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_8_13027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_9_13028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_10_13029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_11_13030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_12_13031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_13_13032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_14_13033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_15_13034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_16_13035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3_13036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_4_13037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_5_13038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_6_13039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_7_13040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_8_13041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_9_13042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_10_13043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_11_13044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_12_13045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_13_13046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_14_13047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_15_13048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_16_13049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3_13050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_4_13051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_5_13052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_6_13053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_7_13054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_8_13055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_9_13056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_10_13057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_11_13058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_12_13059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_13_13060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_14_13061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_15_13062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_16_13063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3_13064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_4_13065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_5_13066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_6_13067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_7_13068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_8_13069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_9_13070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_10_13071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_11_13072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_12_13073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_13_13074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_14_13075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_15_13076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_16_13077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3_13078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_4_13079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_5_13080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_6_13081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_7_13082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_8_13083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_9_13084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_10_13085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_11_13086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_12_13087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_13_13088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_14_13089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_15_13090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_16_13091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3_13092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_4_13093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_5_13094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_6_13095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_7_13096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_8_13097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_9_13098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_10_13099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_11_13100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_12_13101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_13_13102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_14_13103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_15_13104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_16_13105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3_13106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_4_13107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_5_13108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_6_13109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_7_13110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_8_13111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_9_13112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_10_13113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_11_13114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_12_13115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_13_13116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_14_13117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_15_13118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_16_13119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3_13120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_4_13121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_5_13122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_6_13123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_7_13124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_8_13125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_9_13126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_10_13127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_11_13128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_12_13129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_13_13130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_14_13131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_15_13132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_16_13133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3_13134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_4_13135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_5_13136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_6_13137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_7_13138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_8_13139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_9_13140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_10_13141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_11_13142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_12_13143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_13_13144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_14_13145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_15_13146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_16_13147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3_13148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_4_13149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_5_13150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_6_13151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_7_13152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_8_13153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_9_13154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_10_13155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_11_13156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_12_13157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_13_13158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_14_13159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_15_13160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_16_13161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3_13162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_4_13163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_5_13164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_6_13165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_7_13166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_8_13167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_9_13168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_10_13169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_11_13170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_12_13171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_13_13172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_14_13173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_15_13174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_16_13175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3_13176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_4_13177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_5_13178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_6_13179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_7_13180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_8_13181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_9_13182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_10_13183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_11_13184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_12_13185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_13_13186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_14_13187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_15_13188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_16_13189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3_13190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_4_13191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_5_13192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_6_13193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_7_13194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_8_13195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_9_13196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_10_13197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_11_13198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_12_13199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_13_13200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_14_13201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_15_13202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_16_13203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3_13204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_4_13205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_5_13206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_6_13207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_7_13208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_8_13209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_9_13210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_10_13211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_11_13212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_12_13213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_13_13214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_14_13215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_15_13216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_16_13217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3_13218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_4_13219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_5_13220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_6_13221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_7_13222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_8_13223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_9_13224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_10_13225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_11_13226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_12_13227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_13_13228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_14_13229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_15_13230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_16_13231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3_13232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_4_13233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_5_13234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_6_13235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_7_13236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_8_13237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_9_13238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_10_13239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_11_13240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_12_13241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_13_13242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_14_13243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_15_13244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_16_13245 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(wb_adr_i[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(wb_adr_i[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(wb_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(wb_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(wb_adr_i[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(wb_adr_i[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input7 (.I(wb_adr_i[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input8 (.I(wb_adr_i[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 input9 (.I(wb_adr_i[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input10 (.I(wb_adr_i[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(wb_cyc_i),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(wb_dat_i[0]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(wb_dat_i[10]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(wb_dat_i[11]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(wb_dat_i[12]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(wb_dat_i[13]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(wb_dat_i[14]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(wb_dat_i[15]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(wb_dat_i[16]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(wb_dat_i[17]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(wb_dat_i[18]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input22 (.I(wb_dat_i[19]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(wb_dat_i[1]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(wb_dat_i[20]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(wb_dat_i[21]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(wb_dat_i[22]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(wb_dat_i[23]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(wb_dat_i[24]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(wb_dat_i[25]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(wb_dat_i[26]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(wb_dat_i[27]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(wb_dat_i[28]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(wb_dat_i[29]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(wb_dat_i[2]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input35 (.I(wb_dat_i[30]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input36 (.I(wb_dat_i[31]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input37 (.I(wb_dat_i[3]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input38 (.I(wb_dat_i[4]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input39 (.I(wb_dat_i[5]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(wb_dat_i[6]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input41 (.I(wb_dat_i[7]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(wb_dat_i[8]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(wb_dat_i[9]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input44 (.I(wb_rst_i),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(wb_sel_i[0]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(wb_sel_i[1]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(wb_sel_i[2]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(wb_sel_i[3]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(wb_stb_i),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input50 (.I(wb_we_i),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output51 (.I(net51),
    .Z(wb_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output52 (.I(net52),
    .Z(wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output53 (.I(net53),
    .Z(wb_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output54 (.I(net54),
    .Z(wb_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output55 (.I(net55),
    .Z(wb_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output56 (.I(net56),
    .Z(wb_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output57 (.I(net57),
    .Z(wb_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output58 (.I(net58),
    .Z(wb_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output59 (.I(net59),
    .Z(wb_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output60 (.I(net60),
    .Z(wb_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output61 (.I(net61),
    .Z(wb_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output62 (.I(net62),
    .Z(wb_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output63 (.I(net63),
    .Z(wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output64 (.I(net64),
    .Z(wb_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output65 (.I(net65),
    .Z(wb_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output66 (.I(net66),
    .Z(wb_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output67 (.I(net67),
    .Z(wb_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output68 (.I(net68),
    .Z(wb_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output69 (.I(net69),
    .Z(wb_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output70 (.I(net70),
    .Z(wb_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output71 (.I(net71),
    .Z(wb_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output72 (.I(net72),
    .Z(wb_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output73 (.I(net73),
    .Z(wb_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output74 (.I(net74),
    .Z(wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output75 (.I(net75),
    .Z(wb_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output76 (.I(net76),
    .Z(wb_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output77 (.I(net77),
    .Z(wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output78 (.I(net78),
    .Z(wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output79 (.I(net79),
    .Z(wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output80 (.I(net80),
    .Z(wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output81 (.I(net81),
    .Z(wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output82 (.I(net82),
    .Z(wb_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output83 (.I(net83),
    .Z(wb_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire84 (.I(_2253_),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire85 (.I(_2239_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire86 (.I(_2225_),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire87 (.I(_2198_),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire88 (.I(_2184_),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire89 (.I(_2170_),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire90 (.I(_2156_),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 wire92 (.I(_2128_),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire93 (.I(_2100_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire94 (.I(_2087_),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire95 (.I(_2044_),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire96 (.I(_1989_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire97 (.I(_1975_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 wire98 (.I(_1932_),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap100 (.I(_1686_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap102 (.I(_1471_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap104 (.I(_1468_),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire105 (.I(net106),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap106 (.I(_1465_),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap108 (.I(_1462_),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire110 (.I(_1459_),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap112 (.I(_1456_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap114 (.I(_1453_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire115 (.I(net116),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap116 (.I(_1450_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap117 (.I(net122),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap120 (.I(net121),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap121 (.I(_1385_),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap122 (.I(_1385_),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap124 (.I(_2737_),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew125 (.I(net126),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap126 (.I(_2696_),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew127 (.I(net128),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew128 (.I(_2655_),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap130 (.I(_2581_),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap132 (.I(_2540_),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew133 (.I(_2477_),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire134 (.I(_2453_),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew135 (.I(net136),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap136 (.I(_2427_),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire137 (.I(net138),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap138 (.I(_2378_),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew139 (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire141 (.I(_2329_),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire143 (.I(_2274_),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire144 (.I(_2252_),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire145 (.I(_2243_),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire146 (.I(_2218_),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire148 (.I(_2197_),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire150 (.I(_2099_),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire151 (.I(_1936_),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire152 (.I(_1931_),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire153 (.I(_1901_),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire154 (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire155 (.I(_1895_),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire156 (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire157 (.I(_1887_),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire158 (.I(_1864_),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap159 (.I(_1768_),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew160 (.I(net161),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap161 (.I(_1593_),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire162 (.I(net163),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap163 (.I(_1535_),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap164 (.I(net165),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap165 (.I(_1447_),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap166 (.I(_1447_),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew167 (.I(_1384_),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew168 (.I(net169),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap169 (.I(_2512_),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire170 (.I(net171),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire171 (.I(_2476_),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap172 (.I(_2476_),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire173 (.I(net174),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap174 (.I(_2313_),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap176 (.I(_2311_),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap177 (.I(_2284_),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire178 (.I(_2281_),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire179 (.I(_2277_),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire180 (.I(_2270_),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire181 (.I(_2215_),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew182 (.I(net183),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap183 (.I(_1642_),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire184 (.I(_1534_),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap185 (.I(_1477_),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap186 (.I(net187),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap187 (.I(_1390_),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap188 (.I(_1388_),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap189 (.I(\bit_sel[9] ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap190 (.I(\bit_sel[8] ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap191 (.I(\bit_sel[7] ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap192 (.I(\bit_sel[6] ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap193 (.I(\bit_sel[63] ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap194 (.I(\bit_sel[62] ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap195 (.I(\bit_sel[61] ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap196 (.I(\bit_sel[60] ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap197 (.I(\bit_sel[5] ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 max_cap198 (.I(\bit_sel[59] ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap199 (.I(\bit_sel[58] ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap200 (.I(\bit_sel[57] ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap201 (.I(\bit_sel[56] ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap202 (.I(\bit_sel[55] ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap203 (.I(\bit_sel[54] ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap204 (.I(\bit_sel[53] ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap205 (.I(\bit_sel[52] ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 max_cap206 (.I(\bit_sel[51] ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 max_cap207 (.I(\bit_sel[50] ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap208 (.I(\bit_sel[4] ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap209 (.I(\bit_sel[49] ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 max_cap210 (.I(\bit_sel[48] ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap211 (.I(\bit_sel[47] ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap212 (.I(\bit_sel[46] ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap213 (.I(\bit_sel[45] ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap214 (.I(\bit_sel[44] ),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap215 (.I(\bit_sel[43] ),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap216 (.I(\bit_sel[42] ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap217 (.I(\bit_sel[41] ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap218 (.I(\bit_sel[40] ),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap219 (.I(\bit_sel[3] ),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap220 (.I(\bit_sel[39] ),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap221 (.I(\bit_sel[38] ),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap222 (.I(\bit_sel[37] ),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap223 (.I(\bit_sel[36] ),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap224 (.I(\bit_sel[35] ),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap225 (.I(\bit_sel[34] ),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap226 (.I(\bit_sel[33] ),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap227 (.I(\bit_sel[32] ),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap228 (.I(\bit_sel[31] ),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap229 (.I(\bit_sel[30] ),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap230 (.I(\bit_sel[2] ),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap231 (.I(\bit_sel[29] ),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap232 (.I(\bit_sel[28] ),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap233 (.I(\bit_sel[27] ),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap234 (.I(\bit_sel[26] ),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap235 (.I(\bit_sel[25] ),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap236 (.I(\bit_sel[24] ),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap237 (.I(\bit_sel[23] ),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap238 (.I(\bit_sel[22] ),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap239 (.I(\bit_sel[21] ),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap240 (.I(\bit_sel[20] ),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap241 (.I(\bit_sel[1] ),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap242 (.I(\bit_sel[19] ),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap243 (.I(\bit_sel[18] ),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap244 (.I(\bit_sel[17] ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap245 (.I(\bit_sel[16] ),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap246 (.I(\bit_sel[15] ),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap247 (.I(\bit_sel[14] ),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap248 (.I(\bit_sel[13] ),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap249 (.I(\bit_sel[12] ),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap250 (.I(\bit_sel[11] ),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap251 (.I(\bit_sel[10] ),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap252 (.I(\bit_sel[0] ),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 wire253 (.I(net254),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap254 (.I(_2622_),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap255 (.I(net256),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire256 (.I(_2287_),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire257 (.I(_2280_),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap258 (.I(net259),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap259 (.I(_1675_),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire260 (.I(_1590_),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 max_cap261 (.I(net263),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap262 (.I(net263),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap263 (.I(net267),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire264 (.I(net266),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap265 (.I(net266),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap266 (.I(net366),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap267 (.I(_1589_),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew268 (.I(_1565_),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire269 (.I(_1533_),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire270 (.I(net271),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 wire271 (.I(_1531_),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap272 (.I(net273),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap273 (.I(net274),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap274 (.I(net363),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire275 (.I(net277),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap276 (.I(net277),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap277 (.I(net362),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew278 (.I(net280),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap279 (.I(net280),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire280 (.I(net281),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap281 (.I(_1335_),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 load_slew282 (.I(\state[3] ),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap283 (.I(net284),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire284 (.I(net285),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire285 (.I(\state[1] ),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap286 (.I(net287),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire287 (.I(_1518_),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire288 (.I(_1518_),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire289 (.I(_1493_),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire290 (.I(_1493_),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire291 (.I(_1490_),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire292 (.I(_1490_),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire293 (.I(_1487_),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire294 (.I(_1487_),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew295 (.I(_1484_),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire296 (.I(_1484_),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire297 (.I(_1481_),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire298 (.I(_1481_),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire299 (.I(_1478_),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire300 (.I(_1478_),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap301 (.I(net302),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire302 (.I(net303),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap303 (.I(_1472_),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire304 (.I(net306),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap305 (.I(net306),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire306 (.I(_1443_),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire307 (.I(_1440_),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap308 (.I(_1440_),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire309 (.I(net310),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap310 (.I(_1437_),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire311 (.I(net312),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap312 (.I(_1434_),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire313 (.I(net314),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap314 (.I(_1431_),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire315 (.I(_1428_),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap316 (.I(_1428_),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire317 (.I(_1425_),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap318 (.I(_1425_),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire319 (.I(_1422_),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap320 (.I(_1422_),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire321 (.I(net323),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap322 (.I(net323),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire323 (.I(_1419_),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap324 (.I(_1416_),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire325 (.I(_1413_),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire326 (.I(_1413_),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire327 (.I(_1410_),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire328 (.I(_1410_),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire329 (.I(_1407_),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire330 (.I(_1407_),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew331 (.I(_1404_),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire332 (.I(_1404_),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire333 (.I(_1401_),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire334 (.I(_1401_),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire335 (.I(_1398_),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire336 (.I(_1398_),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire337 (.I(_1395_),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire338 (.I(_1395_),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew339 (.I(_1392_),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire340 (.I(_1392_),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire341 (.I(net342),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire342 (.I(net343),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire343 (.I(net344),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 wire344 (.I(net345),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 max_cap345 (.I(net346),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap346 (.I(_1386_),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 load_slew347 (.I(net348),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap348 (.I(_1367_),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 max_cap349 (.I(net350),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire350 (.I(_1367_),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire351 (.I(net352),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew352 (.I(_1365_),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 load_slew353 (.I(net354),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 max_cap354 (.I(_1365_),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap355 (.I(net9),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap356 (.I(net357),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap357 (.I(net358),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire358 (.I(net359),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap359 (.I(net44),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 load_slew360 (.I(net10),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 max_cap361 (.I(net10),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_19_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_21_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_70_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_72_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_75_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_78_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_79_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_80_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_81_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_82_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_83_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_84_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_85_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_leaf_86_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_12 clkload0 (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkload1 (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 clkload2 (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload3 (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkload4 (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkload5 (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload6 (.I(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload7 (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload8 (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload9 (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload10 (.I(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload11 (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload12 (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload13 (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload14 (.I(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload15 (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload16 (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload17 (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload18 (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload19 (.I(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload20 (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload21 (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload22 (.I(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload23 (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload24 (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload25 (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload26 (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload27 (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload28 (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload29 (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload30 (.I(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 clkload31 (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload32 (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload33 (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload34 (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload35 (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload36 (.I(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload37 (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload38 (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload39 (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload40 (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload41 (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload42 (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload43 (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload44 (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload45 (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload46 (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload47 (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload48 (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload49 (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload50 (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload51 (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload52 (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload53 (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload54 (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 clkload55 (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload56 (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload57 (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload58 (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload59 (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload60 (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload61 (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload62 (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload63 (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload64 (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload65 (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload66 (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload67 (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload68 (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload69 (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload70 (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload71 (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload72 (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload73 (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload74 (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload75 (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload76 (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload77 (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload78 (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload79 (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload80 (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload81 (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload82 (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload83 (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer362 (.I(_1530_),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer363 (.I(net362),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer364 (.I(net362),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer365 (.I(net364),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer366 (.I(_1589_),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer367 (.I(net366),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer368 (.I(_1386_),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer369 (.I(net368),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer370 (.I(net368),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 clone371 (.A1(net8),
    .A2(net7),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer372 (.I(_1472_),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer373 (.I(net372),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer374 (.I(net372),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer375 (.I(net372),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_adr_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(wb_adr_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(wb_adr_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(wb_adr_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(wb_adr_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(wb_adr_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(wb_adr_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(wb_adr_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(wb_adr_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_adr_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wb_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(wb_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(wb_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(wb_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(wb_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(wb_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(wb_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(wb_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(wb_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(wb_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(wb_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(wb_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(wb_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(wb_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(wb_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(wb_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(wb_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(wb_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(wb_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(wb_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(wb_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(wb_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(wb_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(wb_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(wb_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(wb_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(wb_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(wb_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(wb_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(wb_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(wb_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(wb_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(wb_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(wb_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(wb_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(wb_sel_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(wb_sel_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(wb_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(wb_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[9].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[99].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[98].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[97].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[96].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[95].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[94].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[93].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[92].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[91].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[90].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[8].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[89].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[88].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[87].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[86].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[85].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[84].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[83].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[82].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[81].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[80].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[7].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[79].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[78].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[77].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[76].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[75].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[74].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[73].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[72].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[71].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[70].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[6].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[69].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[68].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[67].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[66].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[65].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[64].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[63].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[62].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[61].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[60].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[5].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[59].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[58].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[57].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[56].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[55].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[54].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[53].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[52].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[51].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[511].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[510].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[50].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[509].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[508].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[507].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[506].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[505].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[504].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[503].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[502].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[501].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[500].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[4].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[49].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[499].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[498].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[497].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[496].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[495].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[494].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[493].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[492].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[491].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[490].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[48].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[489].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[488].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[487].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[486].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[485].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[484].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[483].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[482].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[481].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[480].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[47].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[479].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[478].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[477].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[476].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[475].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[474].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[473].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[472].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[471].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[470].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[46].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[469].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[468].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[467].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[466].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[465].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[464].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[463].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[462].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[461].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[460].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[45].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[459].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[458].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[457].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[456].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[455].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[454].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[453].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[452].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[451].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[450].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[44].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[449].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[448].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[447].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[446].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[445].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[444].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[443].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[442].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[441].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[440].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[43].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[439].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[438].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[437].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[436].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[435].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[434].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[433].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[432].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[431].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[430].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[42].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[429].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[428].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[427].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[426].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[425].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[424].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[423].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[422].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[421].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[420].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[41].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[419].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[418].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[417].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[416].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[415].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[414].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[413].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[412].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[411].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[410].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[40].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[409].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[408].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[407].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[406].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[405].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[404].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[403].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[402].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[401].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[400].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[3].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[39].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[399].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[398].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[397].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[396].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[395].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[394].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[393].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[392].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[391].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[390].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[38].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[389].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[388].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[387].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[386].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[385].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[384].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[383].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[382].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[381].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[380].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[37].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[379].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[378].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[377].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[376].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[375].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[374].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[373].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[372].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[371].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[370].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[36].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[369].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[368].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[367].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[366].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[365].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[364].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[363].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[362].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[361].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[360].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[35].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[359].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[358].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[357].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[356].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[355].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[354].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[353].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[352].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[351].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[350].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[34].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[349].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[348].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[347].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[346].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[345].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[344].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[343].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[342].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[341].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[340].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[33].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[339].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[338].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[337].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[336].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[335].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[334].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[333].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[332].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[331].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[330].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[32].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[329].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[328].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[327].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[326].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[325].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[324].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[323].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[322].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[321].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[320].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[31].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[319].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[318].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[317].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[316].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[315].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[314].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[313].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[312].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[311].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[310].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[30].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[309].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[308].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[307].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[306].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[305].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[304].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[303].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[302].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[301].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[300].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[2].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[29].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[299].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[298].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[297].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[296].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[295].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[294].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[293].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[292].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[291].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[290].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[28].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[289].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[288].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[287].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[286].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[285].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[284].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[283].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[282].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[281].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[280].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[27].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[279].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[278].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[277].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[276].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[275].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[274].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[273].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[272].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[271].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[270].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[26].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[269].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[268].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[267].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[266].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[265].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[264].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[263].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[262].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[261].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[260].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[25].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[259].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[258].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[257].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[256].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[255].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[254].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[253].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[252].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[251].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[250].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[24].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[249].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[248].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[247].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[246].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[245].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[244].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[243].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[242].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[241].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[240].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[23].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[239].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[238].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[237].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[236].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[235].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[234].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[233].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[232].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[231].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[230].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[22].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[229].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[228].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[227].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[226].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[225].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[224].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[223].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[222].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[221].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[220].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[21].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[219].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[218].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[217].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[216].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[215].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[214].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[213].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[212].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[211].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[210].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[20].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[209].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[208].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[207].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[206].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[205].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[204].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[203].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[202].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[201].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[200].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[1].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[19].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[199].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[198].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[197].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[196].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[195].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[194].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[193].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[192].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[191].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[190].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[18].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[189].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[188].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[187].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[186].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[185].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[184].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[183].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[182].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[181].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[180].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[17].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[179].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[178].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[177].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[176].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[175].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[174].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[173].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[172].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[171].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[170].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[16].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[169].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[168].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[167].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[166].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[165].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[164].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[163].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[162].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[161].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[160].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[15].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[159].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[158].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[157].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[156].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[155].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[154].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[153].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[152].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[151].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[150].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[14].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[149].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[148].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[147].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[146].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[145].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[144].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[143].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[142].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[141].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[140].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[13].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[139].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[138].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[137].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[136].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[135].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[134].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[133].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[132].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[131].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[130].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[12].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[129].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[128].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[127].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[126].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[125].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[124].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[123].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[122].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[121].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[120].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[11].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[119].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[118].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[117].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[116].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[115].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[114].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[113].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[112].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[111].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[110].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[10].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[109].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[108].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[107].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[106].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[105].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[104].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[103].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[102].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[101].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[100].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[0].prog_disable_keep_cell_S  (.I(write_enable_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__ZN (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap281_I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__C (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__ZN (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap354_I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew352_I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__B (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__B (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__ZN (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__ZN (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire350_I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap348_I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__ZN (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A4 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__ZN (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__ZN (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__Z (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew167_I (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__Z (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap122_I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap121_I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__B (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__ZN (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A3 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A3 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__ZN (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap187_I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__B2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__ZN (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__ZN (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire340_I (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew339_I (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__Z (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire338_I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire337_I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__Z (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire332_I (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew331_I (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__Z (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire330_I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire329_I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__Z (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire328_I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire327_I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__Z (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire326_I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire325_I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__Z (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap324_I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__Z (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap320_I (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire319_I (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__Z (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap318_I (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire317_I (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__Z (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap316_I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire315_I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__Z (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap314_I (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__Z (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap312_I (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__Z (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap310_I (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__Z (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap308_I (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire307_I (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__Z (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap166_I (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap165_I (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__C (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__ZN (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__Z (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__Z (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__Z (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__Z (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__Z (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__Z (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__Z (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__Z (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__ZN (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__Z (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap185_I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__ZN (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire300_I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire299_I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__Z (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire298_I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire297_I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__Z (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire296_I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew295_I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__Z (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire294_I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire293_I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__Z (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire292_I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire291_I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__Z (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire290_I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire289_I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__Z (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire288_I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire287_I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__ZN (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__Z (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__ZN (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__B1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__ZN (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__B2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__ZN (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__B2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__ZN (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__B2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__ZN (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__B2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__ZN (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__B2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__ZN (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__B2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__ZN (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__B2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__ZN (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__ZN (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire269_I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__ZN (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire184_I (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__ZN (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap163_I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__ZN (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__B1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__ZN (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew268_I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__B1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__B1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__B1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__B1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__B1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__B2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__Z (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__Z (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__B2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__ZN (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__B2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__ZN (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__B2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__ZN (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__B2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__ZN (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__B2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__ZN (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__ZN (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__B2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__ZN (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire260_I (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__ZN (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__ZN (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__ZN (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap161_I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__ZN (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__B1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__ZN (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__B1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__ZN (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__B1 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__ZN (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__B1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__ZN (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__B1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__ZN (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__B1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__ZN (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__B1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__ZN (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__B1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__ZN (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap183_I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__ZN (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap259_I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__ZN (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__B1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__B1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__B1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__Z (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A3 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A4 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__ZN (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap100_I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__ZN (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap159_I (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A3 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A3 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__Z (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__ZN (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__ZN (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__ZN (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__ZN (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__B2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__ZN (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__ZN (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__ZN (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__ZN (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__B1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__ZN (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__ZN (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__ZN (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__B1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__ZN (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__ZN (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A2 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__ZN (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__ZN (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__B2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__ZN (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__ZN (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__ZN (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__ZN (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire157_I (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__ZN (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__ZN (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A3 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__ZN (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__ZN (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__ZN (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__ZN (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__ZN (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__ZN (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__ZN (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__ZN (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__B (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__Z (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__ZN (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__ZN (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__ZN (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__ZN (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__ZN (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__ZN (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__ZN (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__ZN (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__ZN (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A3 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__ZN (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire97_I (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__ZN (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__ZN (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__ZN (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire96_I (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__ZN (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__ZN (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__B1 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__ZN (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__ZN (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__ZN (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__B1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__ZN (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__ZN (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__ZN (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__B1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__ZN (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__ZN (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__ZN (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__ZN (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__ZN (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__ZN (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__B1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__ZN (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__ZN (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__ZN (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__B1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__ZN (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__ZN (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__ZN (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire94_I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__ZN (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__ZN (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__ZN (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__B1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__ZN (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__ZN (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__ZN (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__B1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__ZN (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__ZN (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__ZN (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__B1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__ZN (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__B2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__ZN (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__ZN (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__B1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__ZN (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__ZN (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__ZN (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__ZN (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__ZN (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__ZN (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__ZN (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire90_I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__ZN (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__ZN (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__ZN (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__ZN (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__ZN (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__ZN (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__ZN (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__ZN (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__B1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__ZN (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__ZN (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__ZN (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__ZN (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__B1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__ZN (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__ZN (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__B1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__ZN (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__ZN (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__ZN (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__ZN (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__B1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__ZN (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__ZN (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__ZN (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__B1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__ZN (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__ZN (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire84_I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__ZN (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__ZN (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__B1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__ZN (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__ZN (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire180_I (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__Z (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__ZN (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__ZN (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire179_I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__ZN (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__ZN (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire257_I (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__ZN (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire178_I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__ZN (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__ZN (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__ZN (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__ZN (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__B1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__ZN (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__B1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__ZN (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__ZN (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__ZN (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__ZN (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap176_I (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__ZN (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap174_I (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__ZN (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__B1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__B1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__ZN (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__B1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__B1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__ZN (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__B1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__B1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__ZN (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__B1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__B1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__ZN (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__B1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__ZN (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__B1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__ZN (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__B1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__B1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__ZN (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__B1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__B1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__ZN (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap138_I (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__ZN (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__B1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__B1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__ZN (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__ZN (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__B1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__B1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__ZN (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__B1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__B1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__ZN (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__B1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__B1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__ZN (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__B1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__B1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__ZN (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__B1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__B1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__ZN (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__B1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__ZN (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap136_I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__ZN (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire134_I (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__B1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__ZN (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__B1 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__B1 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__ZN (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__B1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__B1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__ZN (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__B1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__B1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__ZN (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__B1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__ZN (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__B1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__B1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__ZN (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__B1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__B1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__ZN (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__B1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__B1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__ZN (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap254_I (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__ZN (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap252_I (.I(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[0].bitsel_buf_keep_cell_Z  (.I(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[0]  (.I(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[0]  (.I(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[0]  (.I(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap251_I (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[10].bitsel_buf_keep_cell_Z  (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[10]  (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[10]  (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[10]  (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[10]  (.I(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap250_I (.I(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[11].bitsel_buf_keep_cell_Z  (.I(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[11]  (.I(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[11]  (.I(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[11]  (.I(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap249_I (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[12].bitsel_buf_keep_cell_Z  (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[12]  (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[12]  (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[12]  (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[12]  (.I(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap248_I (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[13].bitsel_buf_keep_cell_Z  (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[13]  (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[13]  (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[13]  (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[13]  (.I(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap247_I (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[14].bitsel_buf_keep_cell_Z  (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[14]  (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[14]  (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[14]  (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[14]  (.I(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap246_I (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[15].bitsel_buf_keep_cell_Z  (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[15]  (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[15]  (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[15]  (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[15]  (.I(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap245_I (.I(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[16].bitsel_buf_keep_cell_Z  (.I(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[16]  (.I(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[16]  (.I(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[16]  (.I(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap244_I (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[17].bitsel_buf_keep_cell_Z  (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[17]  (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[17]  (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[17]  (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[17]  (.I(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap243_I (.I(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[18].bitsel_buf_keep_cell_Z  (.I(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[18]  (.I(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[18]  (.I(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[18]  (.I(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap242_I (.I(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[19].bitsel_buf_keep_cell_Z  (.I(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[19]  (.I(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[19]  (.I(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[19]  (.I(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap241_I (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[1].bitsel_buf_keep_cell_Z  (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[1]  (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[1]  (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[1]  (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[1]  (.I(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap240_I (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[20].bitsel_buf_keep_cell_Z  (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[20]  (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[20]  (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[20]  (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[20]  (.I(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap239_I (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[21].bitsel_buf_keep_cell_Z  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[21]  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[21]  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[21]  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[21]  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[21]  (.I(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap238_I (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[22].bitsel_buf_keep_cell_Z  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[22]  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[22]  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[22]  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[22]  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[22]  (.I(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap237_I (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[23].bitsel_buf_keep_cell_Z  (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[23]  (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[23]  (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[23]  (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[23]  (.I(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap236_I (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[24].bitsel_buf_keep_cell_Z  (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[24]  (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[24]  (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[24]  (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[24]  (.I(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap235_I (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[25].bitsel_buf_keep_cell_Z  (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[25]  (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[25]  (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[25]  (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[25]  (.I(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap234_I (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[26].bitsel_buf_keep_cell_Z  (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[26]  (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[26]  (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[26]  (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[26]  (.I(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap233_I (.I(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[27].bitsel_buf_keep_cell_Z  (.I(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[27]  (.I(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[27]  (.I(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[27]  (.I(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap232_I (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[28].bitsel_buf_keep_cell_Z  (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[28]  (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[28]  (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[28]  (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[28]  (.I(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap231_I (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[29].bitsel_buf_keep_cell_Z  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[29]  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[29]  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[29]  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[29]  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[29]  (.I(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap230_I (.I(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[2].bitsel_buf_keep_cell_Z  (.I(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[2]  (.I(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[2]  (.I(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[2]  (.I(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap229_I (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[30].bitsel_buf_keep_cell_Z  (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[30]  (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[30]  (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[30]  (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[30]  (.I(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap228_I (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[31].bitsel_buf_keep_cell_Z  (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[31]  (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[31]  (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[31]  (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[31]  (.I(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap227_I (.I(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[32].bitsel_buf_keep_cell_Z  (.I(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[32]  (.I(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[32]  (.I(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[32]  (.I(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap226_I (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[33].bitsel_buf_keep_cell_Z  (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[33]  (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[33]  (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[33]  (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[33]  (.I(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap225_I (.I(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[34].bitsel_buf_keep_cell_Z  (.I(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[34]  (.I(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[34]  (.I(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[34]  (.I(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap224_I (.I(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[35].bitsel_buf_keep_cell_Z  (.I(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[35]  (.I(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[35]  (.I(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[35]  (.I(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap223_I (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[36].bitsel_buf_keep_cell_Z  (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[36]  (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[36]  (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[36]  (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[36]  (.I(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap222_I (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[37].bitsel_buf_keep_cell_Z  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[37]  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[37]  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[37]  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[37]  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[37]  (.I(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap221_I (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[38].bitsel_buf_keep_cell_Z  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[38]  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[38]  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[38]  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[38]  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[38]  (.I(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap220_I (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[39].bitsel_buf_keep_cell_Z  (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[39]  (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[39]  (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[39]  (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[39]  (.I(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap219_I (.I(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[3].bitsel_buf_keep_cell_Z  (.I(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[3]  (.I(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[3]  (.I(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[3]  (.I(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap218_I (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[40].bitsel_buf_keep_cell_Z  (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[40]  (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[40]  (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[40]  (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[40]  (.I(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap217_I (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[41].bitsel_buf_keep_cell_Z  (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[41]  (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[41]  (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[41]  (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[41]  (.I(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap216_I (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[42].bitsel_buf_keep_cell_Z  (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[42]  (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[42]  (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[42]  (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[42]  (.I(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap215_I (.I(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[43].bitsel_buf_keep_cell_Z  (.I(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[43]  (.I(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[43]  (.I(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[43]  (.I(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap214_I (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[44].bitsel_buf_keep_cell_Z  (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[44]  (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[44]  (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[44]  (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[44]  (.I(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap213_I (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[45].bitsel_buf_keep_cell_Z  (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[45]  (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[45]  (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[45]  (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[45]  (.I(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap212_I (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[46].bitsel_buf_keep_cell_Z  (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[46]  (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[46]  (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[46]  (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[46]  (.I(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap211_I (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[47].bitsel_buf_keep_cell_Z  (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[47]  (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[47]  (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[47]  (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[47]  (.I(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap210_I (.I(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[48].bitsel_buf_keep_cell_Z  (.I(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[48]  (.I(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[48]  (.I(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[48]  (.I(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap209_I (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[49].bitsel_buf_keep_cell_Z  (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[49]  (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[49]  (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[49]  (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[49]  (.I(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap208_I (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[4].bitsel_buf_keep_cell_Z  (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[4]  (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[4]  (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[4]  (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[4]  (.I(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap207_I (.I(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[50].bitsel_buf_keep_cell_Z  (.I(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[50]  (.I(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[50]  (.I(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[50]  (.I(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap206_I (.I(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[51].bitsel_buf_keep_cell_Z  (.I(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[51]  (.I(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[51]  (.I(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[51]  (.I(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap205_I (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[52].bitsel_buf_keep_cell_Z  (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[52]  (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[52]  (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[52]  (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[52]  (.I(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap204_I (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[53].bitsel_buf_keep_cell_Z  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[53]  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[53]  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[53]  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[53]  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[53]  (.I(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap203_I (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[54].bitsel_buf_keep_cell_Z  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[54]  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[54]  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[54]  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[54]  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[54]  (.I(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap202_I (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[55].bitsel_buf_keep_cell_Z  (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[55]  (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[55]  (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[55]  (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[55]  (.I(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap201_I (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[56].bitsel_buf_keep_cell_Z  (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[56]  (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[56]  (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[56]  (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[56]  (.I(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap200_I (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[57].bitsel_buf_keep_cell_Z  (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[57]  (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[57]  (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[57]  (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[57]  (.I(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap199_I (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[58].bitsel_buf_keep_cell_Z  (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[58]  (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[58]  (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[58]  (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[58]  (.I(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap198_I (.I(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[59].bitsel_buf_keep_cell_Z  (.I(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[59]  (.I(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[59]  (.I(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[59]  (.I(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap197_I (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[5].bitsel_buf_keep_cell_Z  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[5]  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[5]  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[5]  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[5]  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[5]  (.I(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap196_I (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[60].bitsel_buf_keep_cell_Z  (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[60]  (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[60]  (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[60]  (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[60]  (.I(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap195_I (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[61].bitsel_buf_keep_cell_Z  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[61]  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[61]  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[61]  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[61]  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[61]  (.I(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap194_I (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[62].bitsel_buf_keep_cell_Z  (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[62]  (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[62]  (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[62]  (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[62]  (.I(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap193_I (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[63].bitsel_buf_keep_cell_Z  (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[63]  (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[63]  (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[63]  (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[63]  (.I(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap192_I (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[6].bitsel_buf_keep_cell_Z  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[6]  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[6]  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[6]  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[6]  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[6]  (.I(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap191_I (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[7].bitsel_buf_keep_cell_Z  (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[7]  (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[7]  (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[7]  (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[7]  (.I(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap190_I (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[8].bitsel_buf_keep_cell_Z  (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[8]  (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[8]  (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[8]  (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[8]  (.I(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap189_I (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[9].bitsel_buf_keep_cell_Z  (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[9]  (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_BIT_SEL[9]  (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_BIT_SEL[9]  (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_BIT_SEL[9]  (.I(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[24].bitsel_buf_keep_cell_I  (.I(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__Q (.I(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[56].bitsel_buf_keep_cell_I  (.I(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__Q (.I(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[60].bitsel_buf_keep_cell_I  (.I(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__Q (.I(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk3[8].bitsel_buf_keep_cell_I  (.I(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__Q (.I(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[198].prog_disable_keep_cell_Z  (.I(\col_prog_n[198] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[198] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[1].prog_disable_keep_cell_Z  (.I(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[1]  (.I(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[294].prog_disable_keep_cell_Z  (.I(\col_prog_n[294] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[294] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[295].prog_disable_keep_cell_Z  (.I(\col_prog_n[295] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_COL_PROG_N[7]  (.I(\col_prog_n[295] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[2].prog_disable_keep_cell_Z  (.I(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[2]  (.I(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[320].prog_disable_keep_cell_Z  (.I(\col_prog_n[320] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[0]  (.I(\col_prog_n[320] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[321].prog_disable_keep_cell_Z  (.I(\col_prog_n[321] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[1]  (.I(\col_prog_n[321] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[324].prog_disable_keep_cell_Z  (.I(\col_prog_n[324] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[4]  (.I(\col_prog_n[324] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[325].prog_disable_keep_cell_Z  (.I(\col_prog_n[325] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[5]  (.I(\col_prog_n[325] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[326].prog_disable_keep_cell_Z  (.I(\col_prog_n[326] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[326] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[327].prog_disable_keep_cell_Z  (.I(\col_prog_n[327] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_COL_PROG_N[7]  (.I(\col_prog_n[327] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[3].prog_disable_keep_cell_Z  (.I(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[3]  (.I(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[416].prog_disable_keep_cell_Z  (.I(\col_prog_n[416] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[0]  (.I(\col_prog_n[416] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[417].prog_disable_keep_cell_Z  (.I(\col_prog_n[417] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[1]  (.I(\col_prog_n[417] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[418].prog_disable_keep_cell_Z  (.I(\col_prog_n[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[2]  (.I(\col_prog_n[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[419].prog_disable_keep_cell_Z  (.I(\col_prog_n[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[3]  (.I(\col_prog_n[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[420].prog_disable_keep_cell_Z  (.I(\col_prog_n[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[4]  (.I(\col_prog_n[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[421].prog_disable_keep_cell_Z  (.I(\col_prog_n[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[5]  (.I(\col_prog_n[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[422].prog_disable_keep_cell_Z  (.I(\col_prog_n[422] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[422] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[480].prog_disable_keep_cell_Z  (.I(\col_prog_n[480] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[0]  (.I(\col_prog_n[480] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[481].prog_disable_keep_cell_Z  (.I(\col_prog_n[481] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[1]  (.I(\col_prog_n[481] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[482].prog_disable_keep_cell_Z  (.I(\col_prog_n[482] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[2]  (.I(\col_prog_n[482] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[483].prog_disable_keep_cell_Z  (.I(\col_prog_n[483] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[3]  (.I(\col_prog_n[483] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[484].prog_disable_keep_cell_Z  (.I(\col_prog_n[484] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[4]  (.I(\col_prog_n[484] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[485].prog_disable_keep_cell_Z  (.I(\col_prog_n[485] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[5]  (.I(\col_prog_n[485] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[486].prog_disable_keep_cell_Z  (.I(\col_prog_n[486] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[486] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[487].prog_disable_keep_cell_Z  (.I(\col_prog_n[487] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[7]  (.I(\col_prog_n[487] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[4].prog_disable_keep_cell_Z  (.I(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[4]  (.I(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[505].prog_disable_keep_cell_Z  (.I(\col_prog_n[505] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[25]  (.I(\col_prog_n[505] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[507].prog_disable_keep_cell_Z  (.I(\col_prog_n[507] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[27]  (.I(\col_prog_n[507] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[509].prog_disable_keep_cell_Z  (.I(\col_prog_n[509] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[29]  (.I(\col_prog_n[509] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[511].prog_disable_keep_cell_Z  (.I(\col_prog_n[511] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_COL_PROG_N[31]  (.I(\col_prog_n[511] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[5].prog_disable_keep_cell_Z  (.I(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[5]  (.I(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[64].prog_disable_keep_cell_Z  (.I(\col_prog_n[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[2].efuse_array_COL_PROG_N[0]  (.I(\col_prog_n[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[6].prog_disable_keep_cell_Z  (.I(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[6]  (.I(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[7].prog_disable_keep_cell_Z  (.I(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_COL_PROG_N[7]  (.I(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[130].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[130] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__Q (.I(\col_prog_n_reg[130] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__I (.I(\col_prog_n_reg[130] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[256].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[256] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__Q (.I(\col_prog_n_reg[256] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(\col_prog_n_reg[256] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[32].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__Q (.I(\col_prog_n_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A1 (.I(\col_prog_n_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A2 (.I(\col_prog_n_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[33].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__Q (.I(\col_prog_n_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A1 (.I(\col_prog_n_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A2 (.I(\col_prog_n_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[34].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__Q (.I(\col_prog_n_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__A1 (.I(\col_prog_n_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A2 (.I(\col_prog_n_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[35].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__Q (.I(\col_prog_n_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(\col_prog_n_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A2 (.I(\col_prog_n_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[36].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__Q (.I(\col_prog_n_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A1 (.I(\col_prog_n_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(\col_prog_n_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[37].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__Q (.I(\col_prog_n_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(\col_prog_n_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(\col_prog_n_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[38].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__Q (.I(\col_prog_n_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A1 (.I(\col_prog_n_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A2 (.I(\col_prog_n_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[39].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__Q (.I(\col_prog_n_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A1 (.I(\col_prog_n_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A2 (.I(\col_prog_n_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[418].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__Q (.I(\col_prog_n_reg[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(\col_prog_n_reg[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(\col_prog_n_reg[418] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[419].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__Q (.I(\col_prog_n_reg[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(\col_prog_n_reg[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(\col_prog_n_reg[419] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[420].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__Q (.I(\col_prog_n_reg[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(\col_prog_n_reg[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(\col_prog_n_reg[420] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[421].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__Q (.I(\col_prog_n_reg[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(\col_prog_n_reg[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(\col_prog_n_reg[421] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[423].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[423] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__Q (.I(\col_prog_n_reg[423] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(\col_prog_n_reg[423] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(\col_prog_n_reg[423] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[448].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__Q (.I(\col_prog_n_reg[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(\col_prog_n_reg[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(\col_prog_n_reg[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[449].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__Q (.I(\col_prog_n_reg[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(\col_prog_n_reg[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(\col_prog_n_reg[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[450].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__Q (.I(\col_prog_n_reg[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(\col_prog_n_reg[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(\col_prog_n_reg[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[451].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__Q (.I(\col_prog_n_reg[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(\col_prog_n_reg[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(\col_prog_n_reg[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[452].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[452] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__Q (.I(\col_prog_n_reg[452] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(\col_prog_n_reg[452] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(\col_prog_n_reg[452] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[453].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[453] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__Q (.I(\col_prog_n_reg[453] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(\col_prog_n_reg[453] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(\col_prog_n_reg[453] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[454].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__Q (.I(\col_prog_n_reg[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(\col_prog_n_reg[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(\col_prog_n_reg[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[455].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__Q (.I(\col_prog_n_reg[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(\col_prog_n_reg[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(\col_prog_n_reg[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[65].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__Q (.I(\col_prog_n_reg[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A1 (.I(\col_prog_n_reg[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__A2 (.I(\col_prog_n_reg[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[66].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__Q (.I(\col_prog_n_reg[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(\col_prog_n_reg[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A2 (.I(\col_prog_n_reg[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[67].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__Q (.I(\col_prog_n_reg[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A1 (.I(\col_prog_n_reg[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A2 (.I(\col_prog_n_reg[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[68].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__Q (.I(\col_prog_n_reg[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A1 (.I(\col_prog_n_reg[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(\col_prog_n_reg[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[69].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__Q (.I(\col_prog_n_reg[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__A1 (.I(\col_prog_n_reg[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A2 (.I(\col_prog_n_reg[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[70].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__Q (.I(\col_prog_n_reg[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A1 (.I(\col_prog_n_reg[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(\col_prog_n_reg[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[71].prog_disable_keep_cell_I1  (.I(\col_prog_n_reg[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__Q (.I(\col_prog_n_reg[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A1 (.I(\col_prog_n_reg[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A2 (.I(\col_prog_n_reg[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[0]  (.I(\efuse_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(\efuse_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[10]  (.I(\efuse_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(\efuse_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[0]  (.I(\efuse_out[128] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(\efuse_out[128] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[1]  (.I(\efuse_out[129] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(\efuse_out[129] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[12]  (.I(\efuse_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(\efuse_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[2]  (.I(\efuse_out[130] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(\efuse_out[130] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[5]  (.I(\efuse_out[133] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(\efuse_out[133] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[6]  (.I(\efuse_out[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(\efuse_out[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[8]  (.I(\efuse_out[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(\efuse_out[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[9]  (.I(\efuse_out[137] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(\efuse_out[137] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[12]  (.I(\efuse_out[140] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(\efuse_out[140] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[14]  (.I(\efuse_out[142] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(\efuse_out[142] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[17]  (.I(\efuse_out[145] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(\efuse_out[145] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[19]  (.I(\efuse_out[147] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(\efuse_out[147] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[22]  (.I(\efuse_out[150] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A1 (.I(\efuse_out[150] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[23]  (.I(\efuse_out[151] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(\efuse_out[151] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[24]  (.I(\efuse_out[152] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(\efuse_out[152] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[25]  (.I(\efuse_out[153] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(\efuse_out[153] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[26]  (.I(\efuse_out[154] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(\efuse_out[154] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[27]  (.I(\efuse_out[155] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(\efuse_out[155] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[28]  (.I(\efuse_out[156] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(\efuse_out[156] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[29]  (.I(\efuse_out[157] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(\efuse_out[157] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[30]  (.I(\efuse_out[158] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(\efuse_out[158] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_OUT[31]  (.I(\efuse_out[159] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(\efuse_out[159] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[15]  (.I(\efuse_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(\efuse_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[1]  (.I(\efuse_out[161] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__C1 (.I(\efuse_out[161] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[4]  (.I(\efuse_out[164] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__C1 (.I(\efuse_out[164] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[16]  (.I(\efuse_out[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(\efuse_out[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[12]  (.I(\efuse_out[172] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__C1 (.I(\efuse_out[172] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[16]  (.I(\efuse_out[176] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__C1 (.I(\efuse_out[176] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[17]  (.I(\efuse_out[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(\efuse_out[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[23]  (.I(\efuse_out[183] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__C2 (.I(\efuse_out[183] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[24]  (.I(\efuse_out[184] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__C2 (.I(\efuse_out[184] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[25]  (.I(\efuse_out[185] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__C2 (.I(\efuse_out[185] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[26]  (.I(\efuse_out[186] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(\efuse_out[186] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[27]  (.I(\efuse_out[187] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(\efuse_out[187] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[28]  (.I(\efuse_out[188] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__C2 (.I(\efuse_out[188] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[29]  (.I(\efuse_out[189] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(\efuse_out[189] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[18]  (.I(\efuse_out[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(\efuse_out[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[30]  (.I(\efuse_out[190] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(\efuse_out[190] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_OUT[31]  (.I(\efuse_out[191] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(\efuse_out[191] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[19]  (.I(\efuse_out[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(\efuse_out[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[1]  (.I(\efuse_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(\efuse_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_OUT[21]  (.I(\efuse_out[213] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__B2 (.I(\efuse_out[213] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[22]  (.I(\efuse_out[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(\efuse_out[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_OUT[11]  (.I(\efuse_out[235] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__B2 (.I(\efuse_out[235] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_OUT[13]  (.I(\efuse_out[237] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__B2 (.I(\efuse_out[237] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_OUT[15]  (.I(\efuse_out[239] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__B2 (.I(\efuse_out[239] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[23]  (.I(\efuse_out[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A1 (.I(\efuse_out[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[24]  (.I(\efuse_out[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(\efuse_out[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[4]  (.I(\efuse_out[260] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(\efuse_out[260] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[8]  (.I(\efuse_out[264] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(\efuse_out[264] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[9]  (.I(\efuse_out[265] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(\efuse_out[265] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[11]  (.I(\efuse_out[267] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(\efuse_out[267] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[12]  (.I(\efuse_out[268] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(\efuse_out[268] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[13]  (.I(\efuse_out[269] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(\efuse_out[269] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[26]  (.I(\efuse_out[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(\efuse_out[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[15]  (.I(\efuse_out[271] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(\efuse_out[271] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[20]  (.I(\efuse_out[276] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(\efuse_out[276] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[22]  (.I(\efuse_out[278] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(\efuse_out[278] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[27]  (.I(\efuse_out[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(\efuse_out[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_OUT[27]  (.I(\efuse_out[283] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(\efuse_out[283] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[8]  (.I(\efuse_out[296] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__B2 (.I(\efuse_out[296] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[9]  (.I(\efuse_out[297] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__B2 (.I(\efuse_out[297] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[11]  (.I(\efuse_out[299] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__B2 (.I(\efuse_out[299] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[29]  (.I(\efuse_out[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A1 (.I(\efuse_out[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[2]  (.I(\efuse_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(\efuse_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[13]  (.I(\efuse_out[301] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__B2 (.I(\efuse_out[301] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[15]  (.I(\efuse_out[303] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B2 (.I(\efuse_out[303] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[20]  (.I(\efuse_out[308] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B2 (.I(\efuse_out[308] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[22]  (.I(\efuse_out[310] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__C1 (.I(\efuse_out[310] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[26]  (.I(\efuse_out[314] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__C1 (.I(\efuse_out[314] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_OUT[27]  (.I(\efuse_out[315] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__C1 (.I(\efuse_out[315] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_OUT[1]  (.I(\efuse_out[321] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(\efuse_out[321] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_OUT[3]  (.I(\efuse_out[323] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__B2 (.I(\efuse_out[323] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[0]  (.I(\efuse_out[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__B2 (.I(\efuse_out[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[1]  (.I(\efuse_out[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__B2 (.I(\efuse_out[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_OUT[24]  (.I(\efuse_out[344] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A3 (.I(\efuse_out[344] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[2]  (.I(\efuse_out[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__B2 (.I(\efuse_out[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_OUT[1]  (.I(\efuse_out[353] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__B2 (.I(\efuse_out[353] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_OUT[5]  (.I(\efuse_out[357] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__B2 (.I(\efuse_out[357] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[3]  (.I(\efuse_out[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__C1 (.I(\efuse_out[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[4]  (.I(\efuse_out[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__B2 (.I(\efuse_out[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[6]  (.I(\efuse_out[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__B2 (.I(\efuse_out[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[9]  (.I(\efuse_out[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__B2 (.I(\efuse_out[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[10]  (.I(\efuse_out[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__B2 (.I(\efuse_out[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[0]  (.I(\efuse_out[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(\efuse_out[448] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[1]  (.I(\efuse_out[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__B2 (.I(\efuse_out[449] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[12]  (.I(\efuse_out[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__B2 (.I(\efuse_out[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[2]  (.I(\efuse_out[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__C2 (.I(\efuse_out[450] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[3]  (.I(\efuse_out[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__B2 (.I(\efuse_out[451] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[6]  (.I(\efuse_out[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B2 (.I(\efuse_out[454] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[7]  (.I(\efuse_out[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B2 (.I(\efuse_out[455] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[9]  (.I(\efuse_out[457] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__B2 (.I(\efuse_out[457] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[10]  (.I(\efuse_out[458] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B2 (.I(\efuse_out[458] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[14]  (.I(\efuse_out[462] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B2 (.I(\efuse_out[462] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[15]  (.I(\efuse_out[463] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__B2 (.I(\efuse_out[463] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[16]  (.I(\efuse_out[464] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__B2 (.I(\efuse_out[464] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[18]  (.I(\efuse_out[466] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__B2 (.I(\efuse_out[466] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[20]  (.I(\efuse_out[468] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B2 (.I(\efuse_out[468] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[21]  (.I(\efuse_out[469] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B2 (.I(\efuse_out[469] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[22]  (.I(\efuse_out[470] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B2 (.I(\efuse_out[470] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[23]  (.I(\efuse_out[471] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__C2 (.I(\efuse_out[471] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[24]  (.I(\efuse_out[472] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(\efuse_out[472] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[25]  (.I(\efuse_out[473] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B2 (.I(\efuse_out[473] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[26]  (.I(\efuse_out[474] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B2 (.I(\efuse_out[474] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[28]  (.I(\efuse_out[476] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__C2 (.I(\efuse_out[476] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[29]  (.I(\efuse_out[477] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__C2 (.I(\efuse_out[477] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_OUT[31]  (.I(\efuse_out[479] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__B2 (.I(\efuse_out[479] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[15]  (.I(\efuse_out[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B2 (.I(\efuse_out[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[0]  (.I(\efuse_out[480] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B2 (.I(\efuse_out[480] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[1]  (.I(\efuse_out[481] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(\efuse_out[481] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[2]  (.I(\efuse_out[482] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B2 (.I(\efuse_out[482] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[3]  (.I(\efuse_out[483] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(\efuse_out[483] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[6]  (.I(\efuse_out[486] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(\efuse_out[486] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[7]  (.I(\efuse_out[487] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(\efuse_out[487] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[8]  (.I(\efuse_out[488] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__B2 (.I(\efuse_out[488] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[9]  (.I(\efuse_out[489] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(\efuse_out[489] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[16]  (.I(\efuse_out[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B2 (.I(\efuse_out[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[10]  (.I(\efuse_out[490] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(\efuse_out[490] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[11]  (.I(\efuse_out[491] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__B2 (.I(\efuse_out[491] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[13]  (.I(\efuse_out[493] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B2 (.I(\efuse_out[493] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[14]  (.I(\efuse_out[494] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\efuse_out[494] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[16]  (.I(\efuse_out[496] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(\efuse_out[496] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[17]  (.I(\efuse_out[497] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__B2 (.I(\efuse_out[497] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[18]  (.I(\efuse_out[498] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(\efuse_out[498] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[17]  (.I(\efuse_out[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__B2 (.I(\efuse_out[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[4]  (.I(\efuse_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(\efuse_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[20]  (.I(\efuse_out[500] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(\efuse_out[500] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[21]  (.I(\efuse_out[501] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(\efuse_out[501] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[22]  (.I(\efuse_out[502] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(\efuse_out[502] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[23]  (.I(\efuse_out[503] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__B2 (.I(\efuse_out[503] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[24]  (.I(\efuse_out[504] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B2 (.I(\efuse_out[504] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[25]  (.I(\efuse_out[505] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(\efuse_out[505] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[26]  (.I(\efuse_out[506] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(\efuse_out[506] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[28]  (.I(\efuse_out[508] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__B2 (.I(\efuse_out[508] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[29]  (.I(\efuse_out[509] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B2 (.I(\efuse_out[509] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[18]  (.I(\efuse_out[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__B2 (.I(\efuse_out[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_OUT[30]  (.I(\efuse_out[510] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B2 (.I(\efuse_out[510] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[19]  (.I(\efuse_out[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__B2 (.I(\efuse_out[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[22]  (.I(\efuse_out[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B2 (.I(\efuse_out[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[23]  (.I(\efuse_out[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B2 (.I(\efuse_out[55] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[24]  (.I(\efuse_out[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__B2 (.I(\efuse_out[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[26]  (.I(\efuse_out[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__B2 (.I(\efuse_out[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[27]  (.I(\efuse_out[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__B2 (.I(\efuse_out[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_OUT[29]  (.I(\efuse_out[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B2 (.I(\efuse_out[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[6]  (.I(\efuse_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(\efuse_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_OUT[9]  (.I(\efuse_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(\efuse_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_tie_keep_cell_Z (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[9].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[99].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[98].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[97].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[96].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[95].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[94].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[93].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[92].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[91].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[90].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[8].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[89].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[88].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[87].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[86].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[85].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[84].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[83].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[82].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[81].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[80].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[7].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[79].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[78].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[77].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[76].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[75].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[74].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[73].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[72].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[71].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[70].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[6].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[69].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[68].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[67].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[66].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[65].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[64].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[63].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[62].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[61].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[60].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[5].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[59].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[58].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[57].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[56].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[55].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[54].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[53].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[52].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[51].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[511].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[510].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[50].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[509].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[508].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[507].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[506].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[505].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[504].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[503].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[502].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[501].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[500].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[4].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[49].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[499].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[498].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[497].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[496].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[495].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[494].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[493].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[492].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[491].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[490].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[48].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[489].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[488].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[487].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[486].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[485].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[484].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[483].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[482].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[481].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[480].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[47].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[479].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[478].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[477].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[476].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[475].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[474].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[473].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[472].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[471].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[470].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[46].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[469].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[468].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[467].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[466].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[465].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[464].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[463].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[462].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[461].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[460].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[45].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[459].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[458].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[457].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[456].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[455].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[454].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[453].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[452].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[451].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[450].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[44].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[449].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[448].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[447].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[446].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[445].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[444].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[443].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[442].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[441].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[440].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[43].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[439].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[438].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[437].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[436].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[435].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[434].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[433].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[432].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[431].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[430].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[42].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[429].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[428].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[427].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[426].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[425].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[424].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[423].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[422].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[421].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[420].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[41].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[419].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[418].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[417].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[416].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[415].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[414].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[413].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[412].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[411].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[410].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[40].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[409].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[408].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[407].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[406].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[405].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[404].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[403].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[402].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[401].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[400].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[3].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[39].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[399].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[398].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[397].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[396].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[395].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[394].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[393].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[392].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[391].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[390].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[38].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[389].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[388].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[387].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[386].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[385].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[384].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[383].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[382].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[381].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[380].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[37].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[379].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[378].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[377].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[376].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[375].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[374].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[373].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[372].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[371].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[370].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[36].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[369].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[368].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[367].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[366].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[365].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[364].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[363].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[362].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[361].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[360].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[35].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[359].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[358].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[357].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[356].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[355].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[354].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[353].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[352].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[351].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[350].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[34].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[349].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[348].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[347].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[346].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[345].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[344].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[343].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[342].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[341].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[340].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[33].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[339].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[338].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[337].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[336].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[335].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[334].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[333].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[332].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[331].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[330].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[32].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[329].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[328].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[327].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[326].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[325].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[324].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[323].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[322].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[321].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[320].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[31].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[319].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[318].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[317].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[316].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[315].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[314].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[313].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[312].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[311].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[310].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[30].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[309].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[308].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[307].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[306].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[305].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[304].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[303].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[302].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[301].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[300].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[2].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[29].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[299].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[298].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[297].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[296].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[295].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[294].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[293].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[292].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[291].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[290].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[28].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[289].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[288].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[287].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[286].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[285].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[284].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[283].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[282].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[281].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[280].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[27].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[279].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[278].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[277].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[276].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[275].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[274].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[273].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[272].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[271].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[270].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[26].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[269].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[268].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[267].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[266].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[265].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[264].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[263].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[262].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[261].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[260].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[25].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[259].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[258].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[257].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[256].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[255].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[254].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[253].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[252].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[251].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[250].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[24].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[249].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[248].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[247].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[246].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[245].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[244].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[243].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[242].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[241].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[240].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[23].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[239].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[238].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[237].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[236].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[235].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[234].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[233].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[232].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[231].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[230].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[22].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[229].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[228].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[227].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[226].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[225].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[224].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[223].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[222].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[221].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[220].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[21].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[219].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[218].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[217].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[216].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[215].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[214].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[213].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[212].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[211].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[210].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[20].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[209].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[208].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[207].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[206].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[205].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[204].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[203].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[202].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[201].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[200].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[1].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[19].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[199].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[198].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[197].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[196].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[195].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[194].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[193].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[192].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[191].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[190].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[18].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[189].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[188].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[187].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[186].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[185].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[184].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[183].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[182].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[181].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[180].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[17].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[179].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[178].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[177].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[176].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[175].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[174].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[173].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[172].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[171].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[170].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[16].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[169].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[168].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[167].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[166].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[165].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[164].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[163].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[162].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[161].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[160].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[15].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[159].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[158].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[157].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[156].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[155].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[154].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[153].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[152].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[151].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[150].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[14].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[149].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[148].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[147].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[146].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[145].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[144].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[143].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[142].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[141].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[140].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[13].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[139].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[138].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[137].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[136].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[135].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[134].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[133].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[132].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[131].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[130].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[12].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[129].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[128].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[127].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[126].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[125].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[124].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[123].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[122].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[121].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[120].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[11].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[119].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[118].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[117].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[116].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[115].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[114].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[113].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[112].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[111].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[110].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[10].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[109].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[108].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[107].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[106].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[105].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[104].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[103].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[102].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[101].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[100].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk2[0].prog_disable_keep_cell_I0  (.I(one));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[0].preset_buf_keep_cell_Z  (.I(\preset_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[0].efuse_array_PRESET_N  (.I(\preset_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[14].preset_buf_keep_cell_Z  (.I(\preset_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_PRESET_N  (.I(\preset_n[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[15].preset_buf_keep_cell_Z  (.I(\preset_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_PRESET_N  (.I(\preset_n[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[1].preset_buf_keep_cell_Z  (.I(\preset_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[1].efuse_array_PRESET_N  (.I(\preset_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[0].preset_buf_keep_cell_I  (.I(\preset_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__Q (.I(\preset_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B (.I(\preset_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[0].sense_dly_keep_cell_I  (.I(\sense_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__Q (.I(\sense_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__B (.I(\sense_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_genblk4[3].sense_dly_keep_cell_I  (.I(\sense_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__Q (.I(\sense_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__B (.I(\sense_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew282_I (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__Q (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__B (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__Q (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__B (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__Q (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__Q (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__Q (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__Q (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__Q (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__Q (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__Q (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__Q (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__Q (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__Q (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__Q (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__Q (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__Q (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__Q (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__Q (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__Q (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__Q (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__Q (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A2 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__Q (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__Q (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A2 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__Q (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__Q (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__Q (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_Z (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_Z (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_Z (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_Z (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A4 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_Z (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A3 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_Z (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone371_A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_Z (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone371_A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_Z (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap355_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_Z (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__B (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap361_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew360_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_Z (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__B (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__B (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_Z (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_Z (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_Z (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_Z (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_Z (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_Z (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_Z (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_Z (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_Z (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_Z (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_Z (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_Z (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_Z (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_Z (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_Z (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_Z (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_Z (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_Z (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_Z (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_Z (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_Z (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_Z (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap359_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_Z (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_Z (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_Z (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_Z (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_Z (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_Z (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire84_Z (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire85_Z (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire86_Z (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire87_Z (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A2 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire88_Z (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire89_Z (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire90_Z (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire91_Z (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire92_Z (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire91_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire93_Z (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire94_Z (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__B2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire95_Z (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire96_Z (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__B2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire97_Z (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__B2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire98_Z (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire101_Z (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap102_Z (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire103_Z (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap104_Z (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire103_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire105_Z (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap106_Z (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire105_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire107_Z (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap108_Z (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire107_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire109_Z (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire110_Z (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire109_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__B1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire111_Z (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap112_Z (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire113_Z (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap114_Z (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire115_Z (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap116_Z (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire115_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap117_Z (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__C (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap118_Z (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__C (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap119_Z (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__C (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap120_Z (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__C (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap121_Z (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap120_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__C (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap122_Z (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap117_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__C (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew123_Z (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew125_Z (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap126_Z (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew125_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew127_Z (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew128_Z (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew127_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew129_Z (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew131_Z (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap132_Z (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew133_Z (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire134_Z (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__B1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew135_Z (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap136_Z (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew135_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire137_Z (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew139_Z (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap140_Z (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew139_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire141_Z (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire142_Z (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A3 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire143_Z (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire142_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire144_Z (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__B2 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire145_Z (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire146_Z (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire147_Z (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__B2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire148_Z (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire147_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire149_Z (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__B2 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire150_Z (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire151_Z (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire152_Z (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__B1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire153_Z (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire154_Z (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire155_Z (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire154_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire156_Z (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B2 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire157_Z (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire156_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire158_Z (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap159_Z (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew160_Z (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A2 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap161_Z (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew160_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__A2 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire162_Z (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap164_Z (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__C (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap165_Z (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap164_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__C (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap166_Z (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__C (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew167_Z (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew168_Z (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap169_Z (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew168_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire171_Z (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire170_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire173_Z (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap174_Z (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire173_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire175_Z (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap176_Z (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap177_Z (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire178_Z (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire179_Z (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire180_Z (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__B (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew182_Z (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A2 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap183_Z (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew182_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A2 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire184_Z (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__A2 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A2 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A2 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A2 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap185_Z (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__A2 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap186_Z (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap187_Z (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap186_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__A2 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap188_Z (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__B2 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__B2 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap189_Z (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[9]  (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap190_Z (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[8]  (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap191_Z (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[7]  (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap192_Z (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[6]  (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap193_Z (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[63]  (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap194_Z (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[62]  (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap195_Z (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[61]  (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap196_Z (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[60]  (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap197_Z (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[5]  (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap198_Z (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[59]  (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap199_Z (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[58]  (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap200_Z (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[57]  (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap201_Z (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[56]  (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap202_Z (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[55]  (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap203_Z (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[54]  (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap204_Z (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[53]  (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap205_Z (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[52]  (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap206_Z (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[51]  (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap207_Z (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[50]  (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap208_Z (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[4]  (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap209_Z (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[49]  (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap210_Z (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[48]  (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap211_Z (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[47]  (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap212_Z (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[46]  (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap213_Z (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[45]  (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap214_Z (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[44]  (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap215_Z (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[43]  (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap216_Z (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[42]  (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap217_Z (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[41]  (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap218_Z (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[40]  (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap219_Z (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[3]  (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap220_Z (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[39]  (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap221_Z (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[38]  (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap222_Z (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[37]  (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap223_Z (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[36]  (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap224_Z (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[35]  (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap225_Z (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[34]  (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap226_Z (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[33]  (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap227_Z (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[32]  (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap228_Z (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[31]  (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap229_Z (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[30]  (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap230_Z (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[2]  (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap231_Z (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[29]  (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap232_Z (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[28]  (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap233_Z (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[27]  (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap234_Z (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[26]  (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap235_Z (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[25]  (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap236_Z (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[24]  (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap237_Z (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[23]  (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap238_Z (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[22]  (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap239_Z (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[21]  (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap240_Z (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[20]  (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap241_Z (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[1]  (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap242_Z (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[19]  (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap243_Z (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[18]  (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap244_Z (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[17]  (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap245_Z (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[16]  (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap246_Z (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[15]  (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap247_Z (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[14]  (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap248_Z (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[13]  (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap249_Z (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[12]  (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap250_Z (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[11]  (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap251_Z (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[10]  (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap252_Z (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[15].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[14].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[13].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[12].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[11].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[10].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[9].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[8].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[7].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[6].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[5].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[4].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_efuse_gen_depth[3].efuse_array_BIT_SEL[0]  (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire253_Z (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap254_Z (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire253_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap255_Z (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire256_Z (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap255_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire257_Z (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire260_Z (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A2 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap261_Z (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B1 (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap262_Z (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A3 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__C2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__C2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__A3 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__C1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap263_Z (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap262_I (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__C2 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__B1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap261_I (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__C1 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire264_Z (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__C2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__C1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap265_Z (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__C2 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__C1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__C1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A3 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__C1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__B1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__C1 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap266_Z (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire264_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__C2 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap265_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__C1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__B1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap267_Z (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__C1 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__C1 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__C1 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__C1 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap263_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A3 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__C2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__C2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew268_Z (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__B1 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B1 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire269_Z (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire270_Z (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire271_Z (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire270_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap272_Z (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__C1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__B1 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap273_Z (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap272_I (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__C1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A2 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__C1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__C1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B1 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap274_Z (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap273_I (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__C1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A3 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A2 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A2 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A2 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire275_Z (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B1 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap276_Z (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__B1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__B1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A3 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A3 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__B1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__C1 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap277_Z (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__B1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__B1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__B1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire275_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__B1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap276_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__C1 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew278_Z (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__B (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__B (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__C (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__C (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap279_Z (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__B (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__B (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__B (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__B (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__B (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire280_Z (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap279_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__B (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew278_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__C (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap281_Z (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire280_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__C (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__B (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew282_Z (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__I (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap283_Z (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A2 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire284_Z (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap283_I (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire285_Z (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire284_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A1 (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire289_Z (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__A2 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire290_Z (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire291_Z (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A2 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire292_Z (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire293_Z (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire294_Z (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A2 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew295_Z (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__A2 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A1 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A1 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire296_Z (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire297_Z (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__A2 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire298_Z (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire299_Z (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire300_Z (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap301_Z (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__B1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire302_Z (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap301_I (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A3 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A3 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__B1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap303_Z (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire302_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A3 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__B1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire304_Z (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap305_Z (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A2 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire306_Z (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap305_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire304_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire307_Z (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap308_Z (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__A1 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A1 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A1 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A1 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A2 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire309_Z (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap310_Z (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire309_I (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire311_Z (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap312_Z (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire311_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire313_Z (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap314_Z (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire313_I (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire315_Z (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap316_Z (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__A2 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire317_Z (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap318_Z (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire319_Z (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap320_Z (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A2 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire321_Z (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap322_Z (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire323_Z (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire321_I (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap322_I (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap324_Z (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire325_Z (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire326_Z (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire327_Z (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A2 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire328_Z (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire329_Z (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire330_Z (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew331_Z (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire332_Z (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire333_Z (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire334_Z (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire335_Z (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A2 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire336_Z (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire337_Z (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A2 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire338_Z (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew339_Z (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A1 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__A1 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A1 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire340_Z (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire341_Z (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire342_Z (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire341_I (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A3 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire343_Z (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire342_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire344_Z (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire343_I (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap345_Z (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire344_I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A3 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap346_Z (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap345_I (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew347_Z (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__A2 (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A2 (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap348_Z (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew347_I (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__B (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A3 (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A2 (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap349_Z (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__B (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__C (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire350_Z (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap349_I (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__B (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__B (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__C (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__C (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__C (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__C (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__C (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire351_Z (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__B (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew352_Z (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire351_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__B (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew353_Z (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A1 (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap354_Z (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew353_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap355_Z (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__I (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__B (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__C (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap356_Z (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap357_Z (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap356_I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire358_Z (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap357_I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap359_Z (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire358_I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew360_Z (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__B (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap361_Z (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__B2 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__I (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__B (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__B (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__B (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__B (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload7_I (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_Z (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload38_I (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_Z (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload82_I (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_Z (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload72_I (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_Z (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload44_I (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_Z (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload45_I (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_Z (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload61_I (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_Z (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload17_I (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_Z (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload20_I (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__CLK (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_Z (.I(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload12_I (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_Z (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_Z (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0_0_wb_clk_i_Z (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1_0_wb_clk_i_Z (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload0_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_Z (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload1_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_Z (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_Z (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload2_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_Z (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload3_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_Z (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_Z (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload4_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_Z (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkload5_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_Z (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer364_I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer363_I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap277_I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer362_Z (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__B1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__C1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer365_I (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__B1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__B1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer364_Z (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__B1 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__B1 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer365_Z (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__C2 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__C2 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__B1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer367_Z (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer370_I (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer369_I (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer368_Z (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer370_Z (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__B1 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__B1 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__B1 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__B1 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone371_Z (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer375_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer374_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer373_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B1 (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer372_Z (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__B1 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A2 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A2 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A2 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer374_Z (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B1 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__B1 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer375_Z (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_296_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_302_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_308_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_318_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_5062 ();
endmodule
